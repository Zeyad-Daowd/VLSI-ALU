module verilog_multiplier_route (A,
    B,
    result);
 input [31:0] A;
 input [31:0] B;
 output [63:0] result;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;

 sky130_fd_sc_hd__clkinv_8 _05754_ (.A(net57),
    .Y(_00287_));
 sky130_fd_sc_hd__and4_1 _05755_ (.A(net58),
    .B(net59),
    .C(net12),
    .D(net1),
    .X(_00298_));
 sky130_fd_sc_hd__nand4_1 _05756_ (.A(net33),
    .B(net28),
    .C(net44),
    .D(net27),
    .Y(_00309_));
 sky130_fd_sc_hd__a22o_1 _05757_ (.A1(net33),
    .A2(net28),
    .B1(net44),
    .B2(net27),
    .X(_00320_));
 sky130_fd_sc_hd__and2_1 _05758_ (.A(net55),
    .B(net26),
    .X(_00331_));
 sky130_fd_sc_hd__nand3_1 _05759_ (.A(_00309_),
    .B(_00320_),
    .C(_00331_),
    .Y(_00342_));
 sky130_fd_sc_hd__a21o_1 _05760_ (.A1(_00309_),
    .A2(_00320_),
    .B1(_00331_),
    .X(_00353_));
 sky130_fd_sc_hd__and4_1 _05761_ (.A(net33),
    .B(net44),
    .C(net27),
    .D(net26),
    .X(_00364_));
 sky130_fd_sc_hd__nand2_1 _05762_ (.A(net55),
    .B(net23),
    .Y(_00375_));
 sky130_fd_sc_hd__a22oi_2 _05763_ (.A1(net33),
    .A2(net27),
    .B1(net26),
    .B2(net44),
    .Y(_00385_));
 sky130_fd_sc_hd__or3_1 _05764_ (.A(_00364_),
    .B(_00375_),
    .C(_00385_),
    .X(_00396_));
 sky130_fd_sc_hd__o21bai_1 _05765_ (.A1(_00375_),
    .A2(_00385_),
    .B1_N(_00364_),
    .Y(_00407_));
 sky130_fd_sc_hd__and3_1 _05766_ (.A(_00342_),
    .B(_00353_),
    .C(_00407_),
    .X(_00418_));
 sky130_fd_sc_hd__a21o_1 _05767_ (.A1(_00342_),
    .A2(_00353_),
    .B1(_00407_),
    .X(_00429_));
 sky130_fd_sc_hd__nand2b_1 _05768_ (.A_N(_00418_),
    .B(_00429_),
    .Y(_00440_));
 sky130_fd_sc_hd__and4_1 _05769_ (.A(net23),
    .B(net58),
    .C(net59),
    .D(net12),
    .X(_00451_));
 sky130_fd_sc_hd__a22oi_1 _05770_ (.A1(net23),
    .A2(net58),
    .B1(net59),
    .B2(net12),
    .Y(_00462_));
 sky130_fd_sc_hd__or2_1 _05771_ (.A(_00451_),
    .B(_00462_),
    .X(_00473_));
 sky130_fd_sc_hd__nand2_1 _05772_ (.A(net60),
    .B(net1),
    .Y(_00484_));
 sky130_fd_sc_hd__xor2_1 _05773_ (.A(_00473_),
    .B(_00484_),
    .X(_00495_));
 sky130_fd_sc_hd__xor2_1 _05774_ (.A(_00440_),
    .B(_00495_),
    .X(_00505_));
 sky130_fd_sc_hd__o21ai_1 _05775_ (.A1(_00364_),
    .A2(_00385_),
    .B1(_00375_),
    .Y(_00516_));
 sky130_fd_sc_hd__and4_1 _05776_ (.A(net33),
    .B(net44),
    .C(net26),
    .D(net23),
    .X(_00527_));
 sky130_fd_sc_hd__nand2_1 _05777_ (.A(net55),
    .B(net12),
    .Y(_00538_));
 sky130_fd_sc_hd__a22oi_1 _05778_ (.A1(net33),
    .A2(net26),
    .B1(net23),
    .B2(net44),
    .Y(_00549_));
 sky130_fd_sc_hd__nor2_1 _05779_ (.A(_00527_),
    .B(_00549_),
    .Y(_00560_));
 sky130_fd_sc_hd__o21bai_1 _05780_ (.A1(_00538_),
    .A2(_00549_),
    .B1_N(_00527_),
    .Y(_00571_));
 sky130_fd_sc_hd__and3_1 _05781_ (.A(_00396_),
    .B(_00516_),
    .C(_00571_),
    .X(_00582_));
 sky130_fd_sc_hd__a22oi_1 _05782_ (.A1(net58),
    .A2(net12),
    .B1(net1),
    .B2(net59),
    .Y(_00593_));
 sky130_fd_sc_hd__or2_1 _05783_ (.A(_00298_),
    .B(_00593_),
    .X(_00604_));
 sky130_fd_sc_hd__a21oi_1 _05784_ (.A1(_00396_),
    .A2(_00516_),
    .B1(_00571_),
    .Y(_00615_));
 sky130_fd_sc_hd__or3_1 _05785_ (.A(_00582_),
    .B(_00604_),
    .C(_00615_),
    .X(_00626_));
 sky130_fd_sc_hd__nand2b_1 _05786_ (.A_N(_00582_),
    .B(_00626_),
    .Y(_00636_));
 sky130_fd_sc_hd__and2b_1 _05787_ (.A_N(_00505_),
    .B(_00636_),
    .X(_00647_));
 sky130_fd_sc_hd__xnor2_1 _05788_ (.A(_00505_),
    .B(_00636_),
    .Y(_00658_));
 sky130_fd_sc_hd__xnor2_1 _05789_ (.A(_00298_),
    .B(_00658_),
    .Y(_00669_));
 sky130_fd_sc_hd__o21ai_1 _05790_ (.A1(_00582_),
    .A2(_00615_),
    .B1(_00604_),
    .Y(_00680_));
 sky130_fd_sc_hd__and2_1 _05791_ (.A(_00626_),
    .B(_00680_),
    .X(_00691_));
 sky130_fd_sc_hd__xnor2_1 _05792_ (.A(_00538_),
    .B(_00560_),
    .Y(_00702_));
 sky130_fd_sc_hd__and4_1 _05793_ (.A(net33),
    .B(net44),
    .C(net23),
    .D(net12),
    .X(_00713_));
 sky130_fd_sc_hd__a22oi_1 _05794_ (.A1(net33),
    .A2(net23),
    .B1(net12),
    .B2(net44),
    .Y(_00724_));
 sky130_fd_sc_hd__and4bb_1 _05795_ (.A_N(_00713_),
    .B_N(_00724_),
    .C(net55),
    .D(net1),
    .X(_00735_));
 sky130_fd_sc_hd__nor2_1 _05796_ (.A(_00713_),
    .B(_00735_),
    .Y(_00746_));
 sky130_fd_sc_hd__and2b_1 _05797_ (.A_N(_00746_),
    .B(_00702_),
    .X(_00757_));
 sky130_fd_sc_hd__xnor2_1 _05798_ (.A(_00702_),
    .B(_00746_),
    .Y(_00768_));
 sky130_fd_sc_hd__and3_1 _05799_ (.A(net58),
    .B(net1),
    .C(_00768_),
    .X(_00778_));
 sky130_fd_sc_hd__o21ai_1 _05800_ (.A1(_00757_),
    .A2(_00778_),
    .B1(_00691_),
    .Y(_00789_));
 sky130_fd_sc_hd__or3_1 _05801_ (.A(_00691_),
    .B(_00757_),
    .C(_00778_),
    .X(_00800_));
 sky130_fd_sc_hd__a21oi_1 _05802_ (.A1(net58),
    .A2(net1),
    .B1(_00768_),
    .Y(_00811_));
 sky130_fd_sc_hd__nor2_1 _05803_ (.A(_00778_),
    .B(_00811_),
    .Y(_00822_));
 sky130_fd_sc_hd__o2bb2a_1 _05804_ (.A1_N(net55),
    .A2_N(net1),
    .B1(_00713_),
    .B2(_00724_),
    .X(_00833_));
 sky130_fd_sc_hd__nor2_1 _05805_ (.A(_00735_),
    .B(_00833_),
    .Y(_00844_));
 sky130_fd_sc_hd__and2_1 _05806_ (.A(net33),
    .B(net1),
    .X(net65));
 sky130_fd_sc_hd__and3_1 _05807_ (.A(net44),
    .B(net12),
    .C(net65),
    .X(_00865_));
 sky130_fd_sc_hd__and2_1 _05808_ (.A(_00844_),
    .B(_00865_),
    .X(_00876_));
 sky130_fd_sc_hd__and2_1 _05809_ (.A(_00822_),
    .B(_00876_),
    .X(_00887_));
 sky130_fd_sc_hd__nand3_1 _05810_ (.A(_00789_),
    .B(_00800_),
    .C(_00887_),
    .Y(_00898_));
 sky130_fd_sc_hd__or2_1 _05811_ (.A(_00669_),
    .B(_00789_),
    .X(_00909_));
 sky130_fd_sc_hd__nand2_1 _05812_ (.A(_00669_),
    .B(_00789_),
    .Y(_00920_));
 sky130_fd_sc_hd__nand2_1 _05813_ (.A(_00909_),
    .B(_00920_),
    .Y(_00930_));
 sky130_fd_sc_hd__or2_1 _05814_ (.A(_00898_),
    .B(_00930_),
    .X(_00941_));
 sky130_fd_sc_hd__nand2_1 _05815_ (.A(_00898_),
    .B(_00930_),
    .Y(_00952_));
 sky130_fd_sc_hd__and2_1 _05816_ (.A(_00941_),
    .B(_00952_),
    .X(net120));
 sky130_fd_sc_hd__and4_1 _05817_ (.A(net33),
    .B(net28),
    .C(net44),
    .D(net29),
    .X(_00973_));
 sky130_fd_sc_hd__a22oi_2 _05818_ (.A1(net28),
    .A2(net44),
    .B1(net29),
    .B2(net33),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _05819_ (.A(net27),
    .B(net55),
    .Y(_00995_));
 sky130_fd_sc_hd__or3_1 _05820_ (.A(_00973_),
    .B(_00984_),
    .C(_00995_),
    .X(_01006_));
 sky130_fd_sc_hd__o21ai_1 _05821_ (.A1(_00973_),
    .A2(_00984_),
    .B1(_00995_),
    .Y(_01017_));
 sky130_fd_sc_hd__a21bo_1 _05822_ (.A1(_00320_),
    .A2(_00331_),
    .B1_N(_00309_),
    .X(_01028_));
 sky130_fd_sc_hd__nand3_1 _05823_ (.A(_01006_),
    .B(_01017_),
    .C(_01028_),
    .Y(_01039_));
 sky130_fd_sc_hd__a21o_1 _05824_ (.A1(_01006_),
    .A2(_01017_),
    .B1(_01028_),
    .X(_01050_));
 sky130_fd_sc_hd__and4_1 _05825_ (.A(net26),
    .B(net23),
    .C(net58),
    .D(net59),
    .X(_01061_));
 sky130_fd_sc_hd__a22oi_1 _05826_ (.A1(net26),
    .A2(net58),
    .B1(net59),
    .B2(net23),
    .Y(_01071_));
 sky130_fd_sc_hd__nor2_1 _05827_ (.A(_01061_),
    .B(_01071_),
    .Y(_01082_));
 sky130_fd_sc_hd__nand2_1 _05828_ (.A(net12),
    .B(net60),
    .Y(_01093_));
 sky130_fd_sc_hd__xnor2_1 _05829_ (.A(_01082_),
    .B(_01093_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand3_1 _05830_ (.A(_01039_),
    .B(_01050_),
    .C(_01104_),
    .Y(_01115_));
 sky130_fd_sc_hd__a21o_1 _05831_ (.A1(_01039_),
    .A2(_01050_),
    .B1(_01104_),
    .X(_01126_));
 sky130_fd_sc_hd__a21o_1 _05832_ (.A1(_00429_),
    .A2(_00495_),
    .B1(_00418_),
    .X(_01137_));
 sky130_fd_sc_hd__and3_1 _05833_ (.A(_01115_),
    .B(_01126_),
    .C(_01137_),
    .X(_01148_));
 sky130_fd_sc_hd__nand3_1 _05834_ (.A(_01115_),
    .B(_01126_),
    .C(_01137_),
    .Y(_01159_));
 sky130_fd_sc_hd__a21o_1 _05835_ (.A1(_01115_),
    .A2(_01126_),
    .B1(_01137_),
    .X(_01170_));
 sky130_fd_sc_hd__o21bai_1 _05836_ (.A1(_00462_),
    .A2(_00484_),
    .B1_N(_00451_),
    .Y(_01181_));
 sky130_fd_sc_hd__nand2_1 _05837_ (.A(net1),
    .B(net61),
    .Y(_01192_));
 sky130_fd_sc_hd__and3_1 _05838_ (.A(net1),
    .B(net61),
    .C(_01181_),
    .X(_01203_));
 sky130_fd_sc_hd__xnor2_1 _05839_ (.A(_01181_),
    .B(_01192_),
    .Y(_01214_));
 sky130_fd_sc_hd__and3_1 _05840_ (.A(_01159_),
    .B(_01170_),
    .C(_01214_),
    .X(_01224_));
 sky130_fd_sc_hd__a21oi_1 _05841_ (.A1(_01159_),
    .A2(_01170_),
    .B1(_01214_),
    .Y(_01235_));
 sky130_fd_sc_hd__or2_1 _05842_ (.A(_01224_),
    .B(_01235_),
    .X(_01246_));
 sky130_fd_sc_hd__a21oi_1 _05843_ (.A1(_00298_),
    .A2(_00658_),
    .B1(_00647_),
    .Y(_01257_));
 sky130_fd_sc_hd__nor2_1 _05844_ (.A(_01246_),
    .B(_01257_),
    .Y(_01268_));
 sky130_fd_sc_hd__nand2_1 _05845_ (.A(_01246_),
    .B(_01257_),
    .Y(_01279_));
 sky130_fd_sc_hd__nand2b_1 _05846_ (.A_N(_01268_),
    .B(_01279_),
    .Y(_01290_));
 sky130_fd_sc_hd__and3_1 _05847_ (.A(_00909_),
    .B(_00941_),
    .C(_01290_),
    .X(_01301_));
 sky130_fd_sc_hd__a21oi_2 _05848_ (.A1(_00909_),
    .A2(_00941_),
    .B1(_01290_),
    .Y(_01312_));
 sky130_fd_sc_hd__nor2_1 _05849_ (.A(_01301_),
    .B(_01312_),
    .Y(net125));
 sky130_fd_sc_hd__and4_1 _05850_ (.A(net33),
    .B(net44),
    .C(net29),
    .D(net30),
    .X(_01333_));
 sky130_fd_sc_hd__a22oi_2 _05851_ (.A1(net44),
    .A2(net29),
    .B1(net30),
    .B2(net33),
    .Y(_01344_));
 sky130_fd_sc_hd__nand2_1 _05852_ (.A(net28),
    .B(net55),
    .Y(_01355_));
 sky130_fd_sc_hd__or3_1 _05853_ (.A(_01333_),
    .B(_01344_),
    .C(_01355_),
    .X(_01366_));
 sky130_fd_sc_hd__o21ai_1 _05854_ (.A1(_01333_),
    .A2(_01344_),
    .B1(_01355_),
    .Y(_01376_));
 sky130_fd_sc_hd__o21bai_1 _05855_ (.A1(_00984_),
    .A2(_00995_),
    .B1_N(_00973_),
    .Y(_01387_));
 sky130_fd_sc_hd__nand3_1 _05856_ (.A(_01366_),
    .B(_01376_),
    .C(_01387_),
    .Y(_01398_));
 sky130_fd_sc_hd__a21o_1 _05857_ (.A1(_01366_),
    .A2(_01376_),
    .B1(_01387_),
    .X(_01409_));
 sky130_fd_sc_hd__and4_1 _05858_ (.A(net27),
    .B(net26),
    .C(net58),
    .D(net59),
    .X(_01420_));
 sky130_fd_sc_hd__a22o_1 _05859_ (.A1(net27),
    .A2(net58),
    .B1(net59),
    .B2(net26),
    .X(_01431_));
 sky130_fd_sc_hd__and2b_1 _05860_ (.A_N(_01420_),
    .B(_01431_),
    .X(_01442_));
 sky130_fd_sc_hd__nand2_1 _05861_ (.A(net23),
    .B(net60),
    .Y(_01453_));
 sky130_fd_sc_hd__xnor2_1 _05862_ (.A(_01442_),
    .B(_01453_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand3_1 _05863_ (.A(_01398_),
    .B(_01409_),
    .C(_01464_),
    .Y(_01475_));
 sky130_fd_sc_hd__a21o_1 _05864_ (.A1(_01398_),
    .A2(_01409_),
    .B1(_01464_),
    .X(_01486_));
 sky130_fd_sc_hd__a21bo_1 _05865_ (.A1(_01050_),
    .A2(_01104_),
    .B1_N(_01039_),
    .X(_01497_));
 sky130_fd_sc_hd__nand3_2 _05866_ (.A(_01475_),
    .B(_01486_),
    .C(_01497_),
    .Y(_01508_));
 sky130_fd_sc_hd__a21o_1 _05867_ (.A1(_01475_),
    .A2(_01486_),
    .B1(_01497_),
    .X(_01519_));
 sky130_fd_sc_hd__a31o_1 _05868_ (.A1(net12),
    .A2(net60),
    .A3(_01082_),
    .B1(_01061_),
    .X(_01530_));
 sky130_fd_sc_hd__and4_1 _05869_ (.A(net12),
    .B(net1),
    .C(net61),
    .D(net62),
    .X(_01540_));
 sky130_fd_sc_hd__a22oi_1 _05870_ (.A1(net12),
    .A2(net61),
    .B1(net62),
    .B2(net1),
    .Y(_01551_));
 sky130_fd_sc_hd__or2_1 _05871_ (.A(_01540_),
    .B(_01551_),
    .X(_01562_));
 sky130_fd_sc_hd__and2b_1 _05872_ (.A_N(_01562_),
    .B(_01530_),
    .X(_01573_));
 sky130_fd_sc_hd__xnor2_1 _05873_ (.A(_01530_),
    .B(_01562_),
    .Y(_01584_));
 sky130_fd_sc_hd__nand3_2 _05874_ (.A(_01508_),
    .B(_01519_),
    .C(_01584_),
    .Y(_01595_));
 sky130_fd_sc_hd__a21o_1 _05875_ (.A1(_01508_),
    .A2(_01519_),
    .B1(_01584_),
    .X(_01606_));
 sky130_fd_sc_hd__o211ai_4 _05876_ (.A1(_01148_),
    .A2(_01224_),
    .B1(_01595_),
    .C1(_01606_),
    .Y(_01617_));
 sky130_fd_sc_hd__a211o_1 _05877_ (.A1(_01595_),
    .A2(_01606_),
    .B1(_01148_),
    .C1(_01224_),
    .X(_01628_));
 sky130_fd_sc_hd__nand3_2 _05878_ (.A(_01203_),
    .B(_01617_),
    .C(_01628_),
    .Y(_01639_));
 sky130_fd_sc_hd__a21o_1 _05879_ (.A1(_01617_),
    .A2(_01628_),
    .B1(_01203_),
    .X(_01650_));
 sky130_fd_sc_hd__nand3_1 _05880_ (.A(_01268_),
    .B(_01639_),
    .C(_01650_),
    .Y(_01661_));
 sky130_fd_sc_hd__a21o_1 _05881_ (.A1(_01639_),
    .A2(_01650_),
    .B1(_01268_),
    .X(_01672_));
 sky130_fd_sc_hd__nand2_1 _05882_ (.A(_01661_),
    .B(_01672_),
    .Y(_01683_));
 sky130_fd_sc_hd__xnor2_2 _05883_ (.A(_01312_),
    .B(_01683_),
    .Y(net126));
 sky130_fd_sc_hd__or3_1 _05884_ (.A(_00941_),
    .B(_01290_),
    .C(_01683_),
    .X(_01704_));
 sky130_fd_sc_hd__or2_1 _05885_ (.A(_00909_),
    .B(_01290_),
    .X(_01714_));
 sky130_fd_sc_hd__nand2_1 _05886_ (.A(net55),
    .B(net29),
    .Y(_01725_));
 sky130_fd_sc_hd__and4_1 _05887_ (.A(net33),
    .B(net44),
    .C(net30),
    .D(net31),
    .X(_01736_));
 sky130_fd_sc_hd__a22oi_2 _05888_ (.A1(net44),
    .A2(net30),
    .B1(net31),
    .B2(net33),
    .Y(_01747_));
 sky130_fd_sc_hd__or3_1 _05889_ (.A(_01725_),
    .B(_01736_),
    .C(_01747_),
    .X(_01758_));
 sky130_fd_sc_hd__o21ai_1 _05890_ (.A1(_01736_),
    .A2(_01747_),
    .B1(_01725_),
    .Y(_01769_));
 sky130_fd_sc_hd__o21bai_1 _05891_ (.A1(_01344_),
    .A2(_01355_),
    .B1_N(_01333_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand3_1 _05892_ (.A(_01758_),
    .B(_01769_),
    .C(_01780_),
    .Y(_01791_));
 sky130_fd_sc_hd__a21o_1 _05893_ (.A1(_01758_),
    .A2(_01769_),
    .B1(_01780_),
    .X(_01802_));
 sky130_fd_sc_hd__and4_1 _05894_ (.A(net28),
    .B(net27),
    .C(net58),
    .D(net59),
    .X(_01813_));
 sky130_fd_sc_hd__a22oi_1 _05895_ (.A1(net28),
    .A2(net58),
    .B1(net59),
    .B2(net27),
    .Y(_01824_));
 sky130_fd_sc_hd__nor2_1 _05896_ (.A(_01813_),
    .B(_01824_),
    .Y(_01835_));
 sky130_fd_sc_hd__nand2_1 _05897_ (.A(net26),
    .B(net60),
    .Y(_01846_));
 sky130_fd_sc_hd__xnor2_1 _05898_ (.A(_01835_),
    .B(_01846_),
    .Y(_01857_));
 sky130_fd_sc_hd__nand3_1 _05899_ (.A(_01791_),
    .B(_01802_),
    .C(_01857_),
    .Y(_01868_));
 sky130_fd_sc_hd__a21o_1 _05900_ (.A1(_01791_),
    .A2(_01802_),
    .B1(_01857_),
    .X(_01878_));
 sky130_fd_sc_hd__a21bo_1 _05901_ (.A1(_01409_),
    .A2(_01464_),
    .B1_N(_01398_),
    .X(_01889_));
 sky130_fd_sc_hd__and3_1 _05902_ (.A(_01868_),
    .B(_01878_),
    .C(_01889_),
    .X(_01900_));
 sky130_fd_sc_hd__a21oi_1 _05903_ (.A1(_01868_),
    .A2(_01878_),
    .B1(_01889_),
    .Y(_01911_));
 sky130_fd_sc_hd__a31o_1 _05904_ (.A1(net23),
    .A2(net60),
    .A3(_01431_),
    .B1(_01420_),
    .X(_01922_));
 sky130_fd_sc_hd__and4_1 _05905_ (.A(net23),
    .B(net12),
    .C(net61),
    .D(net62),
    .X(_01933_));
 sky130_fd_sc_hd__a22oi_1 _05906_ (.A1(net23),
    .A2(net61),
    .B1(net62),
    .B2(net12),
    .Y(_01944_));
 sky130_fd_sc_hd__nor2_1 _05907_ (.A(_01933_),
    .B(_01944_),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2_1 _05908_ (.A(net1),
    .B(net63),
    .Y(_01966_));
 sky130_fd_sc_hd__xnor2_1 _05909_ (.A(_01955_),
    .B(_01966_),
    .Y(_01977_));
 sky130_fd_sc_hd__and2_1 _05910_ (.A(_01922_),
    .B(_01977_),
    .X(_01988_));
 sky130_fd_sc_hd__xor2_1 _05911_ (.A(_01922_),
    .B(_01977_),
    .X(_01999_));
 sky130_fd_sc_hd__and2_1 _05912_ (.A(_01540_),
    .B(_01999_),
    .X(_02010_));
 sky130_fd_sc_hd__xnor2_1 _05913_ (.A(_01540_),
    .B(_01999_),
    .Y(_02021_));
 sky130_fd_sc_hd__nor3_2 _05914_ (.A(_01900_),
    .B(_01911_),
    .C(_02021_),
    .Y(_02032_));
 sky130_fd_sc_hd__o21a_1 _05915_ (.A1(_01900_),
    .A2(_01911_),
    .B1(_02021_),
    .X(_02043_));
 sky130_fd_sc_hd__a211o_1 _05916_ (.A1(_01508_),
    .A2(_01595_),
    .B1(_02032_),
    .C1(_02043_),
    .X(_02054_));
 sky130_fd_sc_hd__o211ai_2 _05917_ (.A1(_02032_),
    .A2(_02043_),
    .B1(_01508_),
    .C1(_01595_),
    .Y(_02064_));
 sky130_fd_sc_hd__and3_1 _05918_ (.A(_01573_),
    .B(_02054_),
    .C(_02064_),
    .X(_02075_));
 sky130_fd_sc_hd__nand3_1 _05919_ (.A(_01573_),
    .B(_02054_),
    .C(_02064_),
    .Y(_02086_));
 sky130_fd_sc_hd__a21oi_1 _05920_ (.A1(_02054_),
    .A2(_02064_),
    .B1(_01573_),
    .Y(_02097_));
 sky130_fd_sc_hd__a211oi_2 _05921_ (.A1(_01617_),
    .A2(_01639_),
    .B1(_02075_),
    .C1(_02097_),
    .Y(_02108_));
 sky130_fd_sc_hd__o211a_1 _05922_ (.A1(_02075_),
    .A2(_02097_),
    .B1(_01617_),
    .C1(_01639_),
    .X(_02119_));
 sky130_fd_sc_hd__nor3_1 _05923_ (.A(_01661_),
    .B(_02108_),
    .C(_02119_),
    .Y(_02130_));
 sky130_fd_sc_hd__or3_1 _05924_ (.A(_01661_),
    .B(_02108_),
    .C(_02119_),
    .X(_02141_));
 sky130_fd_sc_hd__o21ai_1 _05925_ (.A1(_02108_),
    .A2(_02119_),
    .B1(_01661_),
    .Y(_02152_));
 sky130_fd_sc_hd__and4bb_1 _05926_ (.A_N(_01683_),
    .B_N(_01714_),
    .C(_02141_),
    .D(_02152_),
    .X(_02163_));
 sky130_fd_sc_hd__o2bb2a_1 _05927_ (.A1_N(_02141_),
    .A2_N(_02152_),
    .B1(_01683_),
    .B2(_01714_),
    .X(_02174_));
 sky130_fd_sc_hd__nor2_1 _05928_ (.A(_02163_),
    .B(_02174_),
    .Y(_02185_));
 sky130_fd_sc_hd__or3_1 _05929_ (.A(_01704_),
    .B(_02163_),
    .C(_02174_),
    .X(_02196_));
 sky130_fd_sc_hd__xnor2_2 _05930_ (.A(_01704_),
    .B(_02185_),
    .Y(net127));
 sky130_fd_sc_hd__o211a_1 _05931_ (.A1(_01988_),
    .A2(_02010_),
    .B1(net1),
    .C1(net64),
    .X(_02217_));
 sky130_fd_sc_hd__a211oi_1 _05932_ (.A1(net1),
    .A2(net64),
    .B1(_01988_),
    .C1(_02010_),
    .Y(_02227_));
 sky130_fd_sc_hd__nor2_1 _05933_ (.A(_02217_),
    .B(_02227_),
    .Y(_02238_));
 sky130_fd_sc_hd__o21ba_1 _05934_ (.A1(_01824_),
    .A2(_01846_),
    .B1_N(_01813_),
    .X(_02249_));
 sky130_fd_sc_hd__nand2_1 _05935_ (.A(net12),
    .B(net63),
    .Y(_02260_));
 sky130_fd_sc_hd__and4_1 _05936_ (.A(net26),
    .B(net23),
    .C(net61),
    .D(net62),
    .X(_02271_));
 sky130_fd_sc_hd__a22oi_1 _05937_ (.A1(net26),
    .A2(net61),
    .B1(net62),
    .B2(net23),
    .Y(_02282_));
 sky130_fd_sc_hd__nor2_1 _05938_ (.A(_02271_),
    .B(_02282_),
    .Y(_02293_));
 sky130_fd_sc_hd__xnor2_1 _05939_ (.A(_02260_),
    .B(_02293_),
    .Y(_02304_));
 sky130_fd_sc_hd__nand2b_1 _05940_ (.A_N(_02249_),
    .B(_02304_),
    .Y(_02315_));
 sky130_fd_sc_hd__xnor2_1 _05941_ (.A(_02249_),
    .B(_02304_),
    .Y(_02326_));
 sky130_fd_sc_hd__o21ba_1 _05942_ (.A1(_01944_),
    .A2(_01966_),
    .B1_N(_01933_),
    .X(_02337_));
 sky130_fd_sc_hd__nand2b_1 _05943_ (.A_N(_02337_),
    .B(_02326_),
    .Y(_02348_));
 sky130_fd_sc_hd__xnor2_1 _05944_ (.A(_02326_),
    .B(_02337_),
    .Y(_02359_));
 sky130_fd_sc_hd__and4_1 _05945_ (.A(net28),
    .B(net58),
    .C(net59),
    .D(net29),
    .X(_02370_));
 sky130_fd_sc_hd__a22oi_1 _05946_ (.A1(net28),
    .A2(net59),
    .B1(net29),
    .B2(net58),
    .Y(_02381_));
 sky130_fd_sc_hd__nor2_1 _05947_ (.A(_02370_),
    .B(_02381_),
    .Y(_02392_));
 sky130_fd_sc_hd__nand2_1 _05948_ (.A(net27),
    .B(net60),
    .Y(_02402_));
 sky130_fd_sc_hd__xnor2_1 _05949_ (.A(_02392_),
    .B(_02402_),
    .Y(_02413_));
 sky130_fd_sc_hd__nand2_1 _05950_ (.A(net55),
    .B(net30),
    .Y(_02424_));
 sky130_fd_sc_hd__and4_1 _05951_ (.A(net33),
    .B(net44),
    .C(net31),
    .D(net32),
    .X(_02435_));
 sky130_fd_sc_hd__a22oi_2 _05952_ (.A1(net44),
    .A2(net31),
    .B1(net32),
    .B2(net33),
    .Y(_02446_));
 sky130_fd_sc_hd__or3_1 _05953_ (.A(_02424_),
    .B(_02435_),
    .C(_02446_),
    .X(_02457_));
 sky130_fd_sc_hd__o21ai_1 _05954_ (.A1(_02435_),
    .A2(_02446_),
    .B1(_02424_),
    .Y(_02468_));
 sky130_fd_sc_hd__o21bai_1 _05955_ (.A1(_01725_),
    .A2(_01747_),
    .B1_N(_01736_),
    .Y(_02479_));
 sky130_fd_sc_hd__nand3_1 _05956_ (.A(_02457_),
    .B(_02468_),
    .C(_02479_),
    .Y(_02490_));
 sky130_fd_sc_hd__a21o_1 _05957_ (.A1(_02457_),
    .A2(_02468_),
    .B1(_02479_),
    .X(_02501_));
 sky130_fd_sc_hd__nand3_1 _05958_ (.A(_02413_),
    .B(_02490_),
    .C(_02501_),
    .Y(_02512_));
 sky130_fd_sc_hd__a21o_1 _05959_ (.A1(_02490_),
    .A2(_02501_),
    .B1(_02413_),
    .X(_02523_));
 sky130_fd_sc_hd__a21bo_1 _05960_ (.A1(_01802_),
    .A2(_01857_),
    .B1_N(_01791_),
    .X(_02534_));
 sky130_fd_sc_hd__nand3_2 _05961_ (.A(_02512_),
    .B(_02523_),
    .C(_02534_),
    .Y(_02545_));
 sky130_fd_sc_hd__a21o_1 _05962_ (.A1(_02512_),
    .A2(_02523_),
    .B1(_02534_),
    .X(_02556_));
 sky130_fd_sc_hd__nand3_2 _05963_ (.A(_02359_),
    .B(_02545_),
    .C(_02556_),
    .Y(_02566_));
 sky130_fd_sc_hd__a21o_1 _05964_ (.A1(_02545_),
    .A2(_02556_),
    .B1(_02359_),
    .X(_02577_));
 sky130_fd_sc_hd__o211a_1 _05965_ (.A1(_01900_),
    .A2(_02032_),
    .B1(_02566_),
    .C1(_02577_),
    .X(_02588_));
 sky130_fd_sc_hd__o211ai_1 _05966_ (.A1(_01900_),
    .A2(_02032_),
    .B1(_02566_),
    .C1(_02577_),
    .Y(_02599_));
 sky130_fd_sc_hd__a211o_1 _05967_ (.A1(_02566_),
    .A2(_02577_),
    .B1(_01900_),
    .C1(_02032_),
    .X(_02610_));
 sky130_fd_sc_hd__and3_1 _05968_ (.A(_02238_),
    .B(_02599_),
    .C(_02610_),
    .X(_02621_));
 sky130_fd_sc_hd__a21oi_1 _05969_ (.A1(_02599_),
    .A2(_02610_),
    .B1(_02238_),
    .Y(_02632_));
 sky130_fd_sc_hd__a211o_1 _05970_ (.A1(_02054_),
    .A2(_02086_),
    .B1(_02621_),
    .C1(_02632_),
    .X(_02643_));
 sky130_fd_sc_hd__o211ai_1 _05971_ (.A1(_02621_),
    .A2(_02632_),
    .B1(_02054_),
    .C1(_02086_),
    .Y(_02654_));
 sky130_fd_sc_hd__and3_1 _05972_ (.A(_02108_),
    .B(_02643_),
    .C(_02654_),
    .X(_02665_));
 sky130_fd_sc_hd__inv_2 _05973_ (.A(_02665_),
    .Y(_02676_));
 sky130_fd_sc_hd__a21o_1 _05974_ (.A1(_02643_),
    .A2(_02654_),
    .B1(_02108_),
    .X(_02687_));
 sky130_fd_sc_hd__and2b_1 _05975_ (.A_N(_02665_),
    .B(_02687_),
    .X(_02698_));
 sky130_fd_sc_hd__nand2_1 _05976_ (.A(_02163_),
    .B(_02698_),
    .Y(_02709_));
 sky130_fd_sc_hd__o21ba_1 _05977_ (.A1(_02260_),
    .A2(_02282_),
    .B1_N(_02271_),
    .X(_02720_));
 sky130_fd_sc_hd__o21ba_1 _05978_ (.A1(_02381_),
    .A2(_02402_),
    .B1_N(_02370_),
    .X(_02730_));
 sky130_fd_sc_hd__and4_1 _05979_ (.A(net27),
    .B(net26),
    .C(net61),
    .D(net62),
    .X(_02741_));
 sky130_fd_sc_hd__a22oi_1 _05980_ (.A1(net27),
    .A2(net61),
    .B1(net62),
    .B2(net26),
    .Y(_02752_));
 sky130_fd_sc_hd__nor2_1 _05981_ (.A(_02741_),
    .B(_02752_),
    .Y(_02763_));
 sky130_fd_sc_hd__nand2_1 _05982_ (.A(net23),
    .B(net63),
    .Y(_02774_));
 sky130_fd_sc_hd__xnor2_1 _05983_ (.A(_02763_),
    .B(_02774_),
    .Y(_02785_));
 sky130_fd_sc_hd__nand2b_1 _05984_ (.A_N(_02730_),
    .B(_02785_),
    .Y(_02796_));
 sky130_fd_sc_hd__xnor2_1 _05985_ (.A(_02730_),
    .B(_02785_),
    .Y(_02807_));
 sky130_fd_sc_hd__nand2b_1 _05986_ (.A_N(_02720_),
    .B(_02807_),
    .Y(_02818_));
 sky130_fd_sc_hd__xnor2_1 _05987_ (.A(_02720_),
    .B(_02807_),
    .Y(_02829_));
 sky130_fd_sc_hd__and4_1 _05988_ (.A(net58),
    .B(net59),
    .C(net29),
    .D(net30),
    .X(_02840_));
 sky130_fd_sc_hd__a22oi_1 _05989_ (.A1(net59),
    .A2(net29),
    .B1(net30),
    .B2(net58),
    .Y(_02851_));
 sky130_fd_sc_hd__nor2_1 _05990_ (.A(_02840_),
    .B(_02851_),
    .Y(_02862_));
 sky130_fd_sc_hd__nand2_1 _05991_ (.A(net28),
    .B(net60),
    .Y(_02873_));
 sky130_fd_sc_hd__xnor2_1 _05992_ (.A(_02862_),
    .B(_02873_),
    .Y(_02884_));
 sky130_fd_sc_hd__nand2_1 _05993_ (.A(net55),
    .B(net31),
    .Y(_02894_));
 sky130_fd_sc_hd__and4_1 _05994_ (.A(net33),
    .B(net44),
    .C(net2),
    .D(net32),
    .X(_02905_));
 sky130_fd_sc_hd__a22oi_2 _05995_ (.A1(net33),
    .A2(net2),
    .B1(net32),
    .B2(net44),
    .Y(_02916_));
 sky130_fd_sc_hd__or3_1 _05996_ (.A(_02894_),
    .B(_02905_),
    .C(_02916_),
    .X(_02927_));
 sky130_fd_sc_hd__o21ai_1 _05997_ (.A1(_02905_),
    .A2(_02916_),
    .B1(_02894_),
    .Y(_02938_));
 sky130_fd_sc_hd__o21bai_1 _05998_ (.A1(_02424_),
    .A2(_02446_),
    .B1_N(_02435_),
    .Y(_02949_));
 sky130_fd_sc_hd__nand3_1 _05999_ (.A(_02927_),
    .B(_02938_),
    .C(_02949_),
    .Y(_02960_));
 sky130_fd_sc_hd__a21o_1 _06000_ (.A1(_02927_),
    .A2(_02938_),
    .B1(_02949_),
    .X(_02971_));
 sky130_fd_sc_hd__nand3_1 _06001_ (.A(_02884_),
    .B(_02960_),
    .C(_02971_),
    .Y(_02982_));
 sky130_fd_sc_hd__a21o_1 _06002_ (.A1(_02960_),
    .A2(_02971_),
    .B1(_02884_),
    .X(_02993_));
 sky130_fd_sc_hd__a21bo_1 _06003_ (.A1(_02413_),
    .A2(_02501_),
    .B1_N(_02490_),
    .X(_03004_));
 sky130_fd_sc_hd__nand3_2 _06004_ (.A(_02982_),
    .B(_02993_),
    .C(_03004_),
    .Y(_03015_));
 sky130_fd_sc_hd__a21o_1 _06005_ (.A1(_02982_),
    .A2(_02993_),
    .B1(_03004_),
    .X(_03026_));
 sky130_fd_sc_hd__and3_1 _06006_ (.A(_02829_),
    .B(_03015_),
    .C(_03026_),
    .X(_03037_));
 sky130_fd_sc_hd__nand3_1 _06007_ (.A(_02829_),
    .B(_03015_),
    .C(_03026_),
    .Y(_03047_));
 sky130_fd_sc_hd__a21oi_1 _06008_ (.A1(_03015_),
    .A2(_03026_),
    .B1(_02829_),
    .Y(_03058_));
 sky130_fd_sc_hd__a211o_1 _06009_ (.A1(_02545_),
    .A2(_02566_),
    .B1(_03037_),
    .C1(_03058_),
    .X(_03069_));
 sky130_fd_sc_hd__o211ai_2 _06010_ (.A1(_03037_),
    .A2(_03058_),
    .B1(_02545_),
    .C1(_02566_),
    .Y(_03080_));
 sky130_fd_sc_hd__a22oi_1 _06011_ (.A1(net12),
    .A2(net64),
    .B1(net34),
    .B2(net1),
    .Y(_03091_));
 sky130_fd_sc_hd__and4_1 _06012_ (.A(net12),
    .B(net1),
    .C(net64),
    .D(net34),
    .X(_03102_));
 sky130_fd_sc_hd__or2_1 _06013_ (.A(_03091_),
    .B(_03102_),
    .X(_03113_));
 sky130_fd_sc_hd__a21oi_1 _06014_ (.A1(_02315_),
    .A2(_02348_),
    .B1(_03113_),
    .Y(_03124_));
 sky130_fd_sc_hd__and3_1 _06015_ (.A(_02315_),
    .B(_02348_),
    .C(_03113_),
    .X(_03135_));
 sky130_fd_sc_hd__nor2_1 _06016_ (.A(_03124_),
    .B(_03135_),
    .Y(_03146_));
 sky130_fd_sc_hd__nand3_2 _06017_ (.A(_03069_),
    .B(_03080_),
    .C(_03146_),
    .Y(_03157_));
 sky130_fd_sc_hd__a21o_1 _06018_ (.A1(_03069_),
    .A2(_03080_),
    .B1(_03146_),
    .X(_03168_));
 sky130_fd_sc_hd__o211ai_1 _06019_ (.A1(_02588_),
    .A2(_02621_),
    .B1(_03157_),
    .C1(_03168_),
    .Y(_03179_));
 sky130_fd_sc_hd__a211o_1 _06020_ (.A1(_03157_),
    .A2(_03168_),
    .B1(_02588_),
    .C1(_02621_),
    .X(_03190_));
 sky130_fd_sc_hd__and3_1 _06021_ (.A(_02217_),
    .B(_03179_),
    .C(_03190_),
    .X(_03200_));
 sky130_fd_sc_hd__a21oi_1 _06022_ (.A1(_03179_),
    .A2(_03190_),
    .B1(_02217_),
    .Y(_03211_));
 sky130_fd_sc_hd__or3_2 _06023_ (.A(_02643_),
    .B(_03200_),
    .C(_03211_),
    .X(_03222_));
 sky130_fd_sc_hd__o21ai_2 _06024_ (.A1(_03200_),
    .A2(_03211_),
    .B1(_02643_),
    .Y(_03233_));
 sky130_fd_sc_hd__and2_1 _06025_ (.A(_02130_),
    .B(_02698_),
    .X(_03244_));
 sky130_fd_sc_hd__a21oi_1 _06026_ (.A1(_02130_),
    .A2(_02687_),
    .B1(_02665_),
    .Y(_03255_));
 sky130_fd_sc_hd__nand3_1 _06027_ (.A(_03222_),
    .B(_03233_),
    .C(_03255_),
    .Y(_03266_));
 sky130_fd_sc_hd__a21o_1 _06028_ (.A1(_03222_),
    .A2(_03233_),
    .B1(_03255_),
    .X(_03277_));
 sky130_fd_sc_hd__a21oi_1 _06029_ (.A1(_03266_),
    .A2(_03277_),
    .B1(_02709_),
    .Y(_03288_));
 sky130_fd_sc_hd__a21o_1 _06030_ (.A1(_03266_),
    .A2(_03277_),
    .B1(_02709_),
    .X(_03299_));
 sky130_fd_sc_hd__and3_1 _06031_ (.A(_02709_),
    .B(_03266_),
    .C(_03277_),
    .X(_03310_));
 sky130_fd_sc_hd__nor2_1 _06032_ (.A(_03288_),
    .B(_03310_),
    .Y(_03321_));
 sky130_fd_sc_hd__nor3_1 _06033_ (.A(_02130_),
    .B(_02163_),
    .C(_02698_),
    .Y(_03332_));
 sky130_fd_sc_hd__a211o_1 _06034_ (.A1(_02163_),
    .A2(_02698_),
    .B1(_03244_),
    .C1(_03332_),
    .X(_03343_));
 sky130_fd_sc_hd__nor2_1 _06035_ (.A(_02196_),
    .B(_03343_),
    .Y(_03354_));
 sky130_fd_sc_hd__xor2_2 _06036_ (.A(_03321_),
    .B(_03354_),
    .X(net66));
 sky130_fd_sc_hd__and3_1 _06037_ (.A(_03222_),
    .B(_03233_),
    .C(_03244_),
    .X(_03374_));
 sky130_fd_sc_hd__and4_1 _06038_ (.A(net23),
    .B(net12),
    .C(net64),
    .D(net34),
    .X(_03385_));
 sky130_fd_sc_hd__a22oi_1 _06039_ (.A1(net23),
    .A2(net64),
    .B1(net34),
    .B2(net12),
    .Y(_03396_));
 sky130_fd_sc_hd__nor2_1 _06040_ (.A(_03385_),
    .B(_03396_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2_1 _06041_ (.A(net1),
    .B(net35),
    .Y(_03418_));
 sky130_fd_sc_hd__xnor2_1 _06042_ (.A(_03407_),
    .B(_03418_),
    .Y(_03429_));
 sky130_fd_sc_hd__and2_1 _06043_ (.A(_03102_),
    .B(_03429_),
    .X(_03440_));
 sky130_fd_sc_hd__nor2_1 _06044_ (.A(_03102_),
    .B(_03429_),
    .Y(_03451_));
 sky130_fd_sc_hd__or2_1 _06045_ (.A(_03440_),
    .B(_03451_),
    .X(_03462_));
 sky130_fd_sc_hd__a21oi_1 _06046_ (.A1(_02796_),
    .A2(_02818_),
    .B1(_03462_),
    .Y(_03473_));
 sky130_fd_sc_hd__and3_1 _06047_ (.A(_02796_),
    .B(_02818_),
    .C(_03462_),
    .X(_03484_));
 sky130_fd_sc_hd__nor2_1 _06048_ (.A(_03473_),
    .B(_03484_),
    .Y(_03494_));
 sky130_fd_sc_hd__o21ba_1 _06049_ (.A1(_02752_),
    .A2(_02774_),
    .B1_N(_02741_),
    .X(_03505_));
 sky130_fd_sc_hd__o21ba_1 _06050_ (.A1(_02851_),
    .A2(_02873_),
    .B1_N(_02840_),
    .X(_03516_));
 sky130_fd_sc_hd__and4_1 _06051_ (.A(net28),
    .B(net27),
    .C(net61),
    .D(net62),
    .X(_03527_));
 sky130_fd_sc_hd__a22oi_1 _06052_ (.A1(net28),
    .A2(net61),
    .B1(net62),
    .B2(net27),
    .Y(_03538_));
 sky130_fd_sc_hd__nor2_1 _06053_ (.A(_03527_),
    .B(_03538_),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_1 _06054_ (.A(net26),
    .B(net63),
    .Y(_03560_));
 sky130_fd_sc_hd__xnor2_1 _06055_ (.A(_03549_),
    .B(_03560_),
    .Y(_03571_));
 sky130_fd_sc_hd__nand2b_1 _06056_ (.A_N(_03516_),
    .B(_03571_),
    .Y(_03582_));
 sky130_fd_sc_hd__xnor2_1 _06057_ (.A(_03516_),
    .B(_03571_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2b_1 _06058_ (.A_N(_03505_),
    .B(_03593_),
    .Y(_03604_));
 sky130_fd_sc_hd__xnor2_1 _06059_ (.A(_03505_),
    .B(_03593_),
    .Y(_03615_));
 sky130_fd_sc_hd__nand2_1 _06060_ (.A(net60),
    .B(net29),
    .Y(_03626_));
 sky130_fd_sc_hd__and4_1 _06061_ (.A(net58),
    .B(net59),
    .C(net30),
    .D(net31),
    .X(_03636_));
 sky130_fd_sc_hd__a22oi_1 _06062_ (.A1(net59),
    .A2(net30),
    .B1(net31),
    .B2(net58),
    .Y(_03647_));
 sky130_fd_sc_hd__nor2_1 _06063_ (.A(_03636_),
    .B(_03647_),
    .Y(_03658_));
 sky130_fd_sc_hd__xnor2_1 _06064_ (.A(_03626_),
    .B(_03658_),
    .Y(_03669_));
 sky130_fd_sc_hd__nand2_1 _06065_ (.A(net55),
    .B(net32),
    .Y(_03680_));
 sky130_fd_sc_hd__and4_1 _06066_ (.A(net33),
    .B(net44),
    .C(net2),
    .D(net3),
    .X(_03691_));
 sky130_fd_sc_hd__a22oi_2 _06067_ (.A1(net44),
    .A2(net2),
    .B1(net3),
    .B2(net33),
    .Y(_03702_));
 sky130_fd_sc_hd__or3_1 _06068_ (.A(_03680_),
    .B(_03691_),
    .C(_03702_),
    .X(_03713_));
 sky130_fd_sc_hd__o21ai_1 _06069_ (.A1(_03691_),
    .A2(_03702_),
    .B1(_03680_),
    .Y(_03724_));
 sky130_fd_sc_hd__o21bai_1 _06070_ (.A1(_02894_),
    .A2(_02916_),
    .B1_N(_02905_),
    .Y(_03735_));
 sky130_fd_sc_hd__nand3_1 _06071_ (.A(_03713_),
    .B(_03724_),
    .C(_03735_),
    .Y(_03746_));
 sky130_fd_sc_hd__a21o_1 _06072_ (.A1(_03713_),
    .A2(_03724_),
    .B1(_03735_),
    .X(_03756_));
 sky130_fd_sc_hd__nand3_1 _06073_ (.A(_03669_),
    .B(_03746_),
    .C(_03756_),
    .Y(_03767_));
 sky130_fd_sc_hd__a21o_1 _06074_ (.A1(_03746_),
    .A2(_03756_),
    .B1(_03669_),
    .X(_03778_));
 sky130_fd_sc_hd__a21bo_1 _06075_ (.A1(_02884_),
    .A2(_02971_),
    .B1_N(_02960_),
    .X(_03789_));
 sky130_fd_sc_hd__nand3_1 _06076_ (.A(_03767_),
    .B(_03778_),
    .C(_03789_),
    .Y(_03800_));
 sky130_fd_sc_hd__inv_2 _06077_ (.A(_03800_),
    .Y(_03811_));
 sky130_fd_sc_hd__a21o_1 _06078_ (.A1(_03767_),
    .A2(_03778_),
    .B1(_03789_),
    .X(_03822_));
 sky130_fd_sc_hd__and3_1 _06079_ (.A(_03615_),
    .B(_03800_),
    .C(_03822_),
    .X(_03833_));
 sky130_fd_sc_hd__a21oi_1 _06080_ (.A1(_03800_),
    .A2(_03822_),
    .B1(_03615_),
    .Y(_03844_));
 sky130_fd_sc_hd__a211o_1 _06081_ (.A1(_03015_),
    .A2(_03047_),
    .B1(_03833_),
    .C1(_03844_),
    .X(_03855_));
 sky130_fd_sc_hd__o211ai_2 _06082_ (.A1(_03833_),
    .A2(_03844_),
    .B1(_03015_),
    .C1(_03047_),
    .Y(_03866_));
 sky130_fd_sc_hd__and3_1 _06083_ (.A(_03494_),
    .B(_03855_),
    .C(_03866_),
    .X(_03877_));
 sky130_fd_sc_hd__a21oi_1 _06084_ (.A1(_03855_),
    .A2(_03866_),
    .B1(_03494_),
    .Y(_03887_));
 sky130_fd_sc_hd__a211o_2 _06085_ (.A1(_03069_),
    .A2(_03157_),
    .B1(_03877_),
    .C1(_03887_),
    .X(_03898_));
 sky130_fd_sc_hd__o211ai_2 _06086_ (.A1(_03877_),
    .A2(_03887_),
    .B1(_03069_),
    .C1(_03157_),
    .Y(_03909_));
 sky130_fd_sc_hd__nand3_2 _06087_ (.A(_03124_),
    .B(_03898_),
    .C(_03909_),
    .Y(_03920_));
 sky130_fd_sc_hd__a21o_1 _06088_ (.A1(_03898_),
    .A2(_03909_),
    .B1(_03124_),
    .X(_03931_));
 sky130_fd_sc_hd__and2_1 _06089_ (.A(_03920_),
    .B(_03931_),
    .X(_03942_));
 sky130_fd_sc_hd__a21bo_1 _06090_ (.A1(_02217_),
    .A2(_03190_),
    .B1_N(_03179_),
    .X(_03953_));
 sky130_fd_sc_hd__nand2_1 _06091_ (.A(_03942_),
    .B(_03953_),
    .Y(_03964_));
 sky130_fd_sc_hd__xnor2_1 _06092_ (.A(_03942_),
    .B(_03953_),
    .Y(_03975_));
 sky130_fd_sc_hd__a21boi_1 _06093_ (.A1(_02665_),
    .A2(_03233_),
    .B1_N(_03222_),
    .Y(_03986_));
 sky130_fd_sc_hd__nor2_1 _06094_ (.A(_03222_),
    .B(_03975_),
    .Y(_03997_));
 sky130_fd_sc_hd__and4bb_1 _06095_ (.A_N(_02676_),
    .B_N(_03975_),
    .C(_03233_),
    .D(_03222_),
    .X(_04007_));
 sky130_fd_sc_hd__xnor2_1 _06096_ (.A(_03975_),
    .B(_03986_),
    .Y(_04018_));
 sky130_fd_sc_hd__nand2b_1 _06097_ (.A_N(_04018_),
    .B(_03374_),
    .Y(_04029_));
 sky130_fd_sc_hd__xnor2_2 _06098_ (.A(_03374_),
    .B(_04018_),
    .Y(_04040_));
 sky130_fd_sc_hd__o31ai_2 _06099_ (.A1(_02196_),
    .A2(_03310_),
    .A3(_03343_),
    .B1(_03299_),
    .Y(_04051_));
 sky130_fd_sc_hd__xor2_2 _06100_ (.A(_04040_),
    .B(_04051_),
    .X(net67));
 sky130_fd_sc_hd__nand2_1 _06101_ (.A(_03582_),
    .B(_03604_),
    .Y(_04072_));
 sky130_fd_sc_hd__and4_1 _06102_ (.A(net26),
    .B(net23),
    .C(net64),
    .D(net34),
    .X(_04083_));
 sky130_fd_sc_hd__a22oi_1 _06103_ (.A1(net26),
    .A2(net64),
    .B1(net34),
    .B2(net23),
    .Y(_04094_));
 sky130_fd_sc_hd__nor2_1 _06104_ (.A(_04083_),
    .B(_04094_),
    .Y(_04105_));
 sky130_fd_sc_hd__nand2_1 _06105_ (.A(net12),
    .B(net35),
    .Y(_04115_));
 sky130_fd_sc_hd__xnor2_1 _06106_ (.A(_04105_),
    .B(_04115_),
    .Y(_04126_));
 sky130_fd_sc_hd__o21ba_1 _06107_ (.A1(_03396_),
    .A2(_03418_),
    .B1_N(_03385_),
    .X(_04137_));
 sky130_fd_sc_hd__nand2b_1 _06108_ (.A_N(_04137_),
    .B(_04126_),
    .Y(_04148_));
 sky130_fd_sc_hd__xnor2_1 _06109_ (.A(_04126_),
    .B(_04137_),
    .Y(_04159_));
 sky130_fd_sc_hd__nand3_2 _06110_ (.A(net1),
    .B(net36),
    .C(_04159_),
    .Y(_04170_));
 sky130_fd_sc_hd__a21o_1 _06111_ (.A1(net1),
    .A2(net36),
    .B1(_04159_),
    .X(_04181_));
 sky130_fd_sc_hd__nand2_1 _06112_ (.A(_04170_),
    .B(_04181_),
    .Y(_04192_));
 sky130_fd_sc_hd__xnor2_1 _06113_ (.A(_04072_),
    .B(_04192_),
    .Y(_04203_));
 sky130_fd_sc_hd__xnor2_1 _06114_ (.A(_03440_),
    .B(_04203_),
    .Y(_04214_));
 sky130_fd_sc_hd__o21ba_1 _06115_ (.A1(_03538_),
    .A2(_03560_),
    .B1_N(_03527_),
    .X(_04224_));
 sky130_fd_sc_hd__o21ba_1 _06116_ (.A1(_03626_),
    .A2(_03647_),
    .B1_N(_03636_),
    .X(_04235_));
 sky130_fd_sc_hd__and4_1 _06117_ (.A(net28),
    .B(net29),
    .C(net61),
    .D(net62),
    .X(_04246_));
 sky130_fd_sc_hd__a22oi_1 _06118_ (.A1(net29),
    .A2(net61),
    .B1(net62),
    .B2(net28),
    .Y(_04257_));
 sky130_fd_sc_hd__nor2_1 _06119_ (.A(_04246_),
    .B(_04257_),
    .Y(_04268_));
 sky130_fd_sc_hd__nand2_1 _06120_ (.A(net27),
    .B(net63),
    .Y(_04279_));
 sky130_fd_sc_hd__xnor2_1 _06121_ (.A(_04268_),
    .B(_04279_),
    .Y(_04290_));
 sky130_fd_sc_hd__and2b_1 _06122_ (.A_N(_04235_),
    .B(_04290_),
    .X(_04301_));
 sky130_fd_sc_hd__xnor2_1 _06123_ (.A(_04235_),
    .B(_04290_),
    .Y(_04312_));
 sky130_fd_sc_hd__and2b_1 _06124_ (.A_N(_04224_),
    .B(_04312_),
    .X(_04323_));
 sky130_fd_sc_hd__xnor2_1 _06125_ (.A(_04224_),
    .B(_04312_),
    .Y(_04334_));
 sky130_fd_sc_hd__nand2_1 _06126_ (.A(net60),
    .B(net30),
    .Y(_04344_));
 sky130_fd_sc_hd__and4_1 _06127_ (.A(net58),
    .B(net59),
    .C(net31),
    .D(net32),
    .X(_04355_));
 sky130_fd_sc_hd__a22oi_1 _06128_ (.A1(net59),
    .A2(net31),
    .B1(net32),
    .B2(net58),
    .Y(_04366_));
 sky130_fd_sc_hd__nor2_1 _06129_ (.A(_04355_),
    .B(_04366_),
    .Y(_04377_));
 sky130_fd_sc_hd__xnor2_1 _06130_ (.A(_04344_),
    .B(_04377_),
    .Y(_04388_));
 sky130_fd_sc_hd__nand2_1 _06131_ (.A(net55),
    .B(net2),
    .Y(_04399_));
 sky130_fd_sc_hd__and4_1 _06132_ (.A(net33),
    .B(net44),
    .C(net3),
    .D(net4),
    .X(_04410_));
 sky130_fd_sc_hd__a22oi_2 _06133_ (.A1(net44),
    .A2(net3),
    .B1(net4),
    .B2(net33),
    .Y(_04421_));
 sky130_fd_sc_hd__or3_1 _06134_ (.A(_04399_),
    .B(_04410_),
    .C(_04421_),
    .X(_04432_));
 sky130_fd_sc_hd__o21ai_1 _06135_ (.A1(_04410_),
    .A2(_04421_),
    .B1(_04399_),
    .Y(_04442_));
 sky130_fd_sc_hd__o21bai_1 _06136_ (.A1(_03680_),
    .A2(_03702_),
    .B1_N(_03691_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand3_1 _06137_ (.A(_04432_),
    .B(_04442_),
    .C(_04453_),
    .Y(_04464_));
 sky130_fd_sc_hd__a21o_1 _06138_ (.A1(_04432_),
    .A2(_04442_),
    .B1(_04453_),
    .X(_04475_));
 sky130_fd_sc_hd__nand3_1 _06139_ (.A(_04388_),
    .B(_04464_),
    .C(_04475_),
    .Y(_04486_));
 sky130_fd_sc_hd__a21o_1 _06140_ (.A1(_04464_),
    .A2(_04475_),
    .B1(_04388_),
    .X(_04497_));
 sky130_fd_sc_hd__a21bo_1 _06141_ (.A1(_03669_),
    .A2(_03756_),
    .B1_N(_03746_),
    .X(_04508_));
 sky130_fd_sc_hd__nand3_2 _06142_ (.A(_04486_),
    .B(_04497_),
    .C(_04508_),
    .Y(_04519_));
 sky130_fd_sc_hd__a21o_1 _06143_ (.A1(_04486_),
    .A2(_04497_),
    .B1(_04508_),
    .X(_04530_));
 sky130_fd_sc_hd__nand3_1 _06144_ (.A(_04334_),
    .B(_04519_),
    .C(_04530_),
    .Y(_04540_));
 sky130_fd_sc_hd__a21o_1 _06145_ (.A1(_04519_),
    .A2(_04530_),
    .B1(_04334_),
    .X(_04551_));
 sky130_fd_sc_hd__o211a_1 _06146_ (.A1(_03811_),
    .A2(_03833_),
    .B1(_04540_),
    .C1(_04551_),
    .X(_04562_));
 sky130_fd_sc_hd__a211oi_1 _06147_ (.A1(_04540_),
    .A2(_04551_),
    .B1(_03811_),
    .C1(_03833_),
    .Y(_04573_));
 sky130_fd_sc_hd__nor2_1 _06148_ (.A(_04562_),
    .B(_04573_),
    .Y(_04584_));
 sky130_fd_sc_hd__xnor2_1 _06149_ (.A(_04214_),
    .B(_04584_),
    .Y(_04595_));
 sky130_fd_sc_hd__a21bo_1 _06150_ (.A1(_03494_),
    .A2(_03866_),
    .B1_N(_03855_),
    .X(_04606_));
 sky130_fd_sc_hd__and2_1 _06151_ (.A(_04595_),
    .B(_04606_),
    .X(_04617_));
 sky130_fd_sc_hd__xor2_1 _06152_ (.A(_04595_),
    .B(_04606_),
    .X(_04627_));
 sky130_fd_sc_hd__and2_1 _06153_ (.A(_03473_),
    .B(_04627_),
    .X(_04638_));
 sky130_fd_sc_hd__nor2_1 _06154_ (.A(_03473_),
    .B(_04627_),
    .Y(_04649_));
 sky130_fd_sc_hd__a211oi_4 _06155_ (.A1(_03898_),
    .A2(_03920_),
    .B1(_04638_),
    .C1(_04649_),
    .Y(_04660_));
 sky130_fd_sc_hd__o211a_1 _06156_ (.A1(_04638_),
    .A2(_04649_),
    .B1(_03898_),
    .C1(_03920_),
    .X(_04671_));
 sky130_fd_sc_hd__or3_4 _06157_ (.A(_03964_),
    .B(_04660_),
    .C(_04671_),
    .X(_04682_));
 sky130_fd_sc_hd__o21ai_2 _06158_ (.A1(_04660_),
    .A2(_04671_),
    .B1(_03964_),
    .Y(_04693_));
 sky130_fd_sc_hd__nand3_4 _06159_ (.A(_03997_),
    .B(_04682_),
    .C(_04693_),
    .Y(_04704_));
 sky130_fd_sc_hd__a21o_1 _06160_ (.A1(_04682_),
    .A2(_04693_),
    .B1(_03997_),
    .X(_04715_));
 sky130_fd_sc_hd__and3_1 _06161_ (.A(_04007_),
    .B(_04704_),
    .C(_04715_),
    .X(_04725_));
 sky130_fd_sc_hd__a21o_1 _06162_ (.A1(_04704_),
    .A2(_04715_),
    .B1(_04007_),
    .X(_04736_));
 sky130_fd_sc_hd__nand2b_1 _06163_ (.A_N(_04725_),
    .B(_04736_),
    .Y(_04747_));
 sky130_fd_sc_hd__a21bo_1 _06164_ (.A1(_04040_),
    .A2(_04051_),
    .B1_N(_04029_),
    .X(_04758_));
 sky130_fd_sc_hd__xnor2_2 _06165_ (.A(_04747_),
    .B(_04758_),
    .Y(net68));
 sky130_fd_sc_hd__a21oi_2 _06166_ (.A1(_04736_),
    .A2(_04758_),
    .B1(_04725_),
    .Y(_04779_));
 sky130_fd_sc_hd__a32oi_2 _06167_ (.A1(_04072_),
    .A2(_04170_),
    .A3(_04181_),
    .B1(_04203_),
    .B2(_03440_),
    .Y(_04790_));
 sky130_fd_sc_hd__a22oi_1 _06168_ (.A1(net12),
    .A2(net36),
    .B1(net37),
    .B2(net1),
    .Y(_04801_));
 sky130_fd_sc_hd__and4_1 _06169_ (.A(net12),
    .B(net1),
    .C(net36),
    .D(net37),
    .X(_04811_));
 sky130_fd_sc_hd__or2_1 _06170_ (.A(_04801_),
    .B(_04811_),
    .X(_04822_));
 sky130_fd_sc_hd__and4_1 _06171_ (.A(net27),
    .B(net26),
    .C(net64),
    .D(net34),
    .X(_04833_));
 sky130_fd_sc_hd__a22oi_1 _06172_ (.A1(net27),
    .A2(net64),
    .B1(net34),
    .B2(net26),
    .Y(_04844_));
 sky130_fd_sc_hd__nor2_1 _06173_ (.A(_04833_),
    .B(_04844_),
    .Y(_04855_));
 sky130_fd_sc_hd__nand2_1 _06174_ (.A(net23),
    .B(net35),
    .Y(_04866_));
 sky130_fd_sc_hd__xnor2_1 _06175_ (.A(_04855_),
    .B(_04866_),
    .Y(_04877_));
 sky130_fd_sc_hd__o21ba_1 _06176_ (.A1(_04094_),
    .A2(_04115_),
    .B1_N(_04083_),
    .X(_04888_));
 sky130_fd_sc_hd__nand2b_1 _06177_ (.A_N(_04888_),
    .B(_04877_),
    .Y(_04898_));
 sky130_fd_sc_hd__xnor2_1 _06178_ (.A(_04877_),
    .B(_04888_),
    .Y(_04909_));
 sky130_fd_sc_hd__nand2b_1 _06179_ (.A_N(_04822_),
    .B(_04909_),
    .Y(_04920_));
 sky130_fd_sc_hd__xnor2_1 _06180_ (.A(_04822_),
    .B(_04909_),
    .Y(_04931_));
 sky130_fd_sc_hd__o21a_1 _06181_ (.A1(_04301_),
    .A2(_04323_),
    .B1(_04931_),
    .X(_04942_));
 sky130_fd_sc_hd__nor3_1 _06182_ (.A(_04301_),
    .B(_04323_),
    .C(_04931_),
    .Y(_04953_));
 sky130_fd_sc_hd__a211oi_2 _06183_ (.A1(_04148_),
    .A2(_04170_),
    .B1(_04942_),
    .C1(_04953_),
    .Y(_04964_));
 sky130_fd_sc_hd__o211a_1 _06184_ (.A1(_04942_),
    .A2(_04953_),
    .B1(_04148_),
    .C1(_04170_),
    .X(_04974_));
 sky130_fd_sc_hd__o21ba_1 _06185_ (.A1(_04257_),
    .A2(_04279_),
    .B1_N(_04246_),
    .X(_04985_));
 sky130_fd_sc_hd__o21ba_1 _06186_ (.A1(_04344_),
    .A2(_04366_),
    .B1_N(_04355_),
    .X(_04996_));
 sky130_fd_sc_hd__and4_1 _06187_ (.A(net29),
    .B(net61),
    .C(net30),
    .D(net62),
    .X(_05007_));
 sky130_fd_sc_hd__a22oi_1 _06188_ (.A1(net61),
    .A2(net30),
    .B1(net62),
    .B2(net29),
    .Y(_05018_));
 sky130_fd_sc_hd__nor2_1 _06189_ (.A(_05007_),
    .B(_05018_),
    .Y(_05029_));
 sky130_fd_sc_hd__nand2_1 _06190_ (.A(net28),
    .B(net63),
    .Y(_05040_));
 sky130_fd_sc_hd__xnor2_1 _06191_ (.A(_05029_),
    .B(_05040_),
    .Y(_05050_));
 sky130_fd_sc_hd__nand2b_1 _06192_ (.A_N(_04996_),
    .B(_05050_),
    .Y(_05061_));
 sky130_fd_sc_hd__xnor2_1 _06193_ (.A(_04996_),
    .B(_05050_),
    .Y(_05072_));
 sky130_fd_sc_hd__nand2b_1 _06194_ (.A_N(_04985_),
    .B(_05072_),
    .Y(_05083_));
 sky130_fd_sc_hd__xnor2_1 _06195_ (.A(_04985_),
    .B(_05072_),
    .Y(_05094_));
 sky130_fd_sc_hd__and4_1 _06196_ (.A(net58),
    .B(net59),
    .C(net2),
    .D(net32),
    .X(_05104_));
 sky130_fd_sc_hd__a22oi_1 _06197_ (.A1(net58),
    .A2(net2),
    .B1(net32),
    .B2(net59),
    .Y(_05115_));
 sky130_fd_sc_hd__nor2_1 _06198_ (.A(_05104_),
    .B(_05115_),
    .Y(_05126_));
 sky130_fd_sc_hd__nand2_1 _06199_ (.A(net60),
    .B(net31),
    .Y(_05137_));
 sky130_fd_sc_hd__xnor2_1 _06200_ (.A(_05126_),
    .B(_05137_),
    .Y(_05148_));
 sky130_fd_sc_hd__nand2_1 _06201_ (.A(net55),
    .B(net3),
    .Y(_05159_));
 sky130_fd_sc_hd__and4_1 _06202_ (.A(net33),
    .B(net44),
    .C(net4),
    .D(net5),
    .X(_05169_));
 sky130_fd_sc_hd__a22oi_2 _06203_ (.A1(net44),
    .A2(net4),
    .B1(net5),
    .B2(net33),
    .Y(_05180_));
 sky130_fd_sc_hd__or3_1 _06204_ (.A(_05159_),
    .B(_05169_),
    .C(_05180_),
    .X(_05191_));
 sky130_fd_sc_hd__o21ai_1 _06205_ (.A1(_05169_),
    .A2(_05180_),
    .B1(_05159_),
    .Y(_05202_));
 sky130_fd_sc_hd__o21bai_1 _06206_ (.A1(_04399_),
    .A2(_04421_),
    .B1_N(_04410_),
    .Y(_05212_));
 sky130_fd_sc_hd__nand3_1 _06207_ (.A(_05191_),
    .B(_05202_),
    .C(_05212_),
    .Y(_05223_));
 sky130_fd_sc_hd__a21o_1 _06208_ (.A1(_05191_),
    .A2(_05202_),
    .B1(_05212_),
    .X(_05234_));
 sky130_fd_sc_hd__nand3_1 _06209_ (.A(_05148_),
    .B(_05223_),
    .C(_05234_),
    .Y(_05245_));
 sky130_fd_sc_hd__a21o_1 _06210_ (.A1(_05223_),
    .A2(_05234_),
    .B1(_05148_),
    .X(_05256_));
 sky130_fd_sc_hd__a21bo_1 _06211_ (.A1(_04388_),
    .A2(_04475_),
    .B1_N(_04464_),
    .X(_05266_));
 sky130_fd_sc_hd__nand3_2 _06212_ (.A(_05245_),
    .B(_05256_),
    .C(_05266_),
    .Y(_05277_));
 sky130_fd_sc_hd__a21o_1 _06213_ (.A1(_05245_),
    .A2(_05256_),
    .B1(_05266_),
    .X(_05288_));
 sky130_fd_sc_hd__and3_1 _06214_ (.A(_05094_),
    .B(_05277_),
    .C(_05288_),
    .X(_05299_));
 sky130_fd_sc_hd__nand3_1 _06215_ (.A(_05094_),
    .B(_05277_),
    .C(_05288_),
    .Y(_05309_));
 sky130_fd_sc_hd__a21oi_1 _06216_ (.A1(_05277_),
    .A2(_05288_),
    .B1(_05094_),
    .Y(_05320_));
 sky130_fd_sc_hd__a211o_1 _06217_ (.A1(_04519_),
    .A2(_04540_),
    .B1(_05299_),
    .C1(_05320_),
    .X(_05331_));
 sky130_fd_sc_hd__o211ai_1 _06218_ (.A1(_05299_),
    .A2(_05320_),
    .B1(_04519_),
    .C1(_04540_),
    .Y(_05341_));
 sky130_fd_sc_hd__or4bb_2 _06219_ (.A(_04964_),
    .B(_04974_),
    .C_N(_05331_),
    .D_N(_05341_),
    .X(_05350_));
 sky130_fd_sc_hd__a2bb2o_1 _06220_ (.A1_N(_04964_),
    .A2_N(_04974_),
    .B1(_05331_),
    .B2(_05341_),
    .X(_05354_));
 sky130_fd_sc_hd__o21bai_1 _06221_ (.A1(_04214_),
    .A2(_04573_),
    .B1_N(_04562_),
    .Y(_05355_));
 sky130_fd_sc_hd__and3_1 _06222_ (.A(_05350_),
    .B(_05354_),
    .C(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__a21oi_1 _06223_ (.A1(_05350_),
    .A2(_05354_),
    .B1(_05355_),
    .Y(_05357_));
 sky130_fd_sc_hd__nor3_1 _06224_ (.A(_04790_),
    .B(_05356_),
    .C(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__o21a_1 _06225_ (.A1(_05356_),
    .A2(_05357_),
    .B1(_04790_),
    .X(_05359_));
 sky130_fd_sc_hd__a21o_1 _06226_ (.A1(_03473_),
    .A2(_04627_),
    .B1(_04617_),
    .X(_05360_));
 sky130_fd_sc_hd__nor3b_1 _06227_ (.A(_05358_),
    .B(_05359_),
    .C_N(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__inv_2 _06228_ (.A(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__o21ba_1 _06229_ (.A1(_05358_),
    .A2(_05359_),
    .B1_N(_05360_),
    .X(_05363_));
 sky130_fd_sc_hd__nor2_1 _06230_ (.A(_05361_),
    .B(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__nand2_1 _06231_ (.A(_04660_),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__xnor2_2 _06232_ (.A(_04660_),
    .B(_05364_),
    .Y(_05366_));
 sky130_fd_sc_hd__nand3_1 _06233_ (.A(_04682_),
    .B(_04704_),
    .C(_05366_),
    .Y(_05367_));
 sky130_fd_sc_hd__or2_1 _06234_ (.A(_04682_),
    .B(_05366_),
    .X(_05368_));
 sky130_fd_sc_hd__o211ai_2 _06235_ (.A1(_04704_),
    .A2(_05366_),
    .B1(_05367_),
    .C1(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__xor2_1 _06236_ (.A(_04779_),
    .B(_05369_),
    .X(net69));
 sky130_fd_sc_hd__o22ai_1 _06237_ (.A1(_04704_),
    .A2(_05366_),
    .B1(_05369_),
    .B2(_04779_),
    .Y(_05370_));
 sky130_fd_sc_hd__o21ai_2 _06238_ (.A1(_04942_),
    .A2(_04964_),
    .B1(_04811_),
    .Y(_05371_));
 sky130_fd_sc_hd__or3_1 _06239_ (.A(_04811_),
    .B(_04942_),
    .C(_04964_),
    .X(_05372_));
 sky130_fd_sc_hd__and2_1 _06240_ (.A(_05371_),
    .B(_05372_),
    .X(_05373_));
 sky130_fd_sc_hd__nand2_1 _06241_ (.A(_04898_),
    .B(_04920_),
    .Y(_05374_));
 sky130_fd_sc_hd__and4_1 _06242_ (.A(net23),
    .B(net12),
    .C(net36),
    .D(net37),
    .X(_05375_));
 sky130_fd_sc_hd__a22oi_1 _06243_ (.A1(net23),
    .A2(net36),
    .B1(net37),
    .B2(net12),
    .Y(_05376_));
 sky130_fd_sc_hd__nor2_1 _06244_ (.A(_05375_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__nand2_1 _06245_ (.A(net1),
    .B(net38),
    .Y(_05378_));
 sky130_fd_sc_hd__xnor2_1 _06246_ (.A(_05377_),
    .B(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__and4_1 _06247_ (.A(net28),
    .B(net27),
    .C(net64),
    .D(net34),
    .X(_05380_));
 sky130_fd_sc_hd__a22oi_1 _06248_ (.A1(net28),
    .A2(net64),
    .B1(net34),
    .B2(net27),
    .Y(_05381_));
 sky130_fd_sc_hd__nor2_1 _06249_ (.A(_05380_),
    .B(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__nand2_1 _06250_ (.A(net26),
    .B(net35),
    .Y(_05383_));
 sky130_fd_sc_hd__xnor2_1 _06251_ (.A(_05382_),
    .B(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__o21ba_1 _06252_ (.A1(_04844_),
    .A2(_04866_),
    .B1_N(_04833_),
    .X(_05385_));
 sky130_fd_sc_hd__and2b_1 _06253_ (.A_N(_05385_),
    .B(_05384_),
    .X(_05386_));
 sky130_fd_sc_hd__xnor2_1 _06254_ (.A(_05384_),
    .B(_05385_),
    .Y(_05387_));
 sky130_fd_sc_hd__and2_1 _06255_ (.A(_05379_),
    .B(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__xnor2_1 _06256_ (.A(_05379_),
    .B(_05387_),
    .Y(_05389_));
 sky130_fd_sc_hd__a21o_1 _06257_ (.A1(_05061_),
    .A2(_05083_),
    .B1(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__nand3_1 _06258_ (.A(_05061_),
    .B(_05083_),
    .C(_05389_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand3_1 _06259_ (.A(_05374_),
    .B(_05390_),
    .C(_05391_),
    .Y(_05392_));
 sky130_fd_sc_hd__a21o_1 _06260_ (.A1(_05390_),
    .A2(_05391_),
    .B1(_05374_),
    .X(_05393_));
 sky130_fd_sc_hd__o21ba_1 _06261_ (.A1(_05018_),
    .A2(_05040_),
    .B1_N(_05007_),
    .X(_05394_));
 sky130_fd_sc_hd__o21ba_1 _06262_ (.A1(_05115_),
    .A2(_05137_),
    .B1_N(_05104_),
    .X(_05395_));
 sky130_fd_sc_hd__and4_1 _06263_ (.A(net61),
    .B(net30),
    .C(net62),
    .D(net31),
    .X(_05396_));
 sky130_fd_sc_hd__a22oi_1 _06264_ (.A1(net30),
    .A2(net62),
    .B1(net31),
    .B2(net61),
    .Y(_05397_));
 sky130_fd_sc_hd__nor2_1 _06265_ (.A(_05396_),
    .B(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__nand2_1 _06266_ (.A(net29),
    .B(net63),
    .Y(_05399_));
 sky130_fd_sc_hd__xnor2_1 _06267_ (.A(_05398_),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__nand2b_1 _06268_ (.A_N(_05395_),
    .B(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__xnor2_1 _06269_ (.A(_05395_),
    .B(_05400_),
    .Y(_05402_));
 sky130_fd_sc_hd__nand2b_1 _06270_ (.A_N(_05394_),
    .B(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__xnor2_1 _06271_ (.A(_05394_),
    .B(_05402_),
    .Y(_05404_));
 sky130_fd_sc_hd__and4_1 _06272_ (.A(net58),
    .B(net59),
    .C(net2),
    .D(net3),
    .X(_05405_));
 sky130_fd_sc_hd__a22oi_1 _06273_ (.A1(net59),
    .A2(net2),
    .B1(net3),
    .B2(net58),
    .Y(_05406_));
 sky130_fd_sc_hd__nor2_1 _06274_ (.A(_05405_),
    .B(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__nand2_1 _06275_ (.A(net60),
    .B(net32),
    .Y(_05408_));
 sky130_fd_sc_hd__xnor2_1 _06276_ (.A(_05407_),
    .B(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__nand2_1 _06277_ (.A(net55),
    .B(net4),
    .Y(_05410_));
 sky130_fd_sc_hd__and4_1 _06278_ (.A(net33),
    .B(net44),
    .C(net5),
    .D(net6),
    .X(_05411_));
 sky130_fd_sc_hd__a22oi_2 _06279_ (.A1(net44),
    .A2(net5),
    .B1(net6),
    .B2(net33),
    .Y(_05412_));
 sky130_fd_sc_hd__or3_1 _06280_ (.A(_05410_),
    .B(_05411_),
    .C(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__o21ai_1 _06281_ (.A1(_05411_),
    .A2(_05412_),
    .B1(_05410_),
    .Y(_05414_));
 sky130_fd_sc_hd__o21bai_1 _06282_ (.A1(_05159_),
    .A2(_05180_),
    .B1_N(_05169_),
    .Y(_05415_));
 sky130_fd_sc_hd__nand3_1 _06283_ (.A(_05413_),
    .B(_05414_),
    .C(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__a21o_1 _06284_ (.A1(_05413_),
    .A2(_05414_),
    .B1(_05415_),
    .X(_05417_));
 sky130_fd_sc_hd__nand3_1 _06285_ (.A(_05409_),
    .B(_05416_),
    .C(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__a21o_1 _06286_ (.A1(_05416_),
    .A2(_05417_),
    .B1(_05409_),
    .X(_05419_));
 sky130_fd_sc_hd__a21bo_1 _06287_ (.A1(_05148_),
    .A2(_05234_),
    .B1_N(_05223_),
    .X(_05420_));
 sky130_fd_sc_hd__nand3_2 _06288_ (.A(_05418_),
    .B(_05419_),
    .C(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__a21o_1 _06289_ (.A1(_05418_),
    .A2(_05419_),
    .B1(_05420_),
    .X(_05422_));
 sky130_fd_sc_hd__and3_1 _06290_ (.A(_05404_),
    .B(_05421_),
    .C(_05422_),
    .X(_05423_));
 sky130_fd_sc_hd__nand3_1 _06291_ (.A(_05404_),
    .B(_05421_),
    .C(_05422_),
    .Y(_05424_));
 sky130_fd_sc_hd__a21oi_1 _06292_ (.A1(_05421_),
    .A2(_05422_),
    .B1(_05404_),
    .Y(_05425_));
 sky130_fd_sc_hd__a211o_1 _06293_ (.A1(_05277_),
    .A2(_05309_),
    .B1(_05423_),
    .C1(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__o211ai_2 _06294_ (.A1(_05423_),
    .A2(_05425_),
    .B1(_05277_),
    .C1(_05309_),
    .Y(_05427_));
 sky130_fd_sc_hd__and4_1 _06295_ (.A(_05392_),
    .B(_05393_),
    .C(_05426_),
    .D(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__nand4_1 _06296_ (.A(_05392_),
    .B(_05393_),
    .C(_05426_),
    .D(_05427_),
    .Y(_05429_));
 sky130_fd_sc_hd__a22oi_1 _06297_ (.A1(_05392_),
    .A2(_05393_),
    .B1(_05426_),
    .B2(_05427_),
    .Y(_05430_));
 sky130_fd_sc_hd__a211o_1 _06298_ (.A1(_05331_),
    .A2(_05350_),
    .B1(_05428_),
    .C1(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__o211ai_1 _06299_ (.A1(_05428_),
    .A2(_05430_),
    .B1(_05331_),
    .C1(_05350_),
    .Y(_05432_));
 sky130_fd_sc_hd__nand3_1 _06300_ (.A(_05373_),
    .B(_05431_),
    .C(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__a21o_1 _06301_ (.A1(_05431_),
    .A2(_05432_),
    .B1(_05373_),
    .X(_05434_));
 sky130_fd_sc_hd__nand2_1 _06302_ (.A(_05433_),
    .B(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__nor2_1 _06303_ (.A(_05356_),
    .B(_05358_),
    .Y(_05436_));
 sky130_fd_sc_hd__nor2_1 _06304_ (.A(_05435_),
    .B(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__xnor2_1 _06305_ (.A(_05435_),
    .B(_05436_),
    .Y(_05438_));
 sky130_fd_sc_hd__or2_1 _06306_ (.A(_05362_),
    .B(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__nand2_1 _06307_ (.A(_05362_),
    .B(_05438_),
    .Y(_05440_));
 sky130_fd_sc_hd__nand2_1 _06308_ (.A(_05439_),
    .B(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__nor2_1 _06309_ (.A(_05365_),
    .B(_05441_),
    .Y(_05442_));
 sky130_fd_sc_hd__nand2_1 _06310_ (.A(_05365_),
    .B(_05368_),
    .Y(_05443_));
 sky130_fd_sc_hd__xnor2_1 _06311_ (.A(_05441_),
    .B(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__xor2_1 _06312_ (.A(_05370_),
    .B(_05444_),
    .X(net70));
 sky130_fd_sc_hd__a2bb2o_1 _06313_ (.A1_N(_05368_),
    .A2_N(_05441_),
    .B1(_05444_),
    .B2(_05370_),
    .X(_05445_));
 sky130_fd_sc_hd__o21ba_1 _06314_ (.A1(_05376_),
    .A2(_05378_),
    .B1_N(_05375_),
    .X(_05446_));
 sky130_fd_sc_hd__nand2_1 _06315_ (.A(net1),
    .B(net39),
    .Y(_05447_));
 sky130_fd_sc_hd__nor2_1 _06316_ (.A(_05446_),
    .B(_05447_),
    .Y(_05448_));
 sky130_fd_sc_hd__xnor2_1 _06317_ (.A(_05446_),
    .B(_05447_),
    .Y(_05449_));
 sky130_fd_sc_hd__a21oi_1 _06318_ (.A1(_05390_),
    .A2(_05392_),
    .B1(_05449_),
    .Y(_05450_));
 sky130_fd_sc_hd__and3_1 _06319_ (.A(_05390_),
    .B(_05392_),
    .C(_05449_),
    .X(_05451_));
 sky130_fd_sc_hd__nor2_1 _06320_ (.A(_05450_),
    .B(_05451_),
    .Y(_05452_));
 sky130_fd_sc_hd__and4_1 _06321_ (.A(net26),
    .B(net23),
    .C(net36),
    .D(net37),
    .X(_05453_));
 sky130_fd_sc_hd__a22oi_1 _06322_ (.A1(net26),
    .A2(net36),
    .B1(net37),
    .B2(net23),
    .Y(_05454_));
 sky130_fd_sc_hd__nor2_1 _06323_ (.A(_05453_),
    .B(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__a21oi_1 _06324_ (.A1(net12),
    .A2(net38),
    .B1(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__and3_1 _06325_ (.A(net12),
    .B(net38),
    .C(_05455_),
    .X(_05457_));
 sky130_fd_sc_hd__nor2_1 _06326_ (.A(_05456_),
    .B(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__and4_1 _06327_ (.A(net28),
    .B(net29),
    .C(net64),
    .D(net34),
    .X(_05459_));
 sky130_fd_sc_hd__a22o_1 _06328_ (.A1(net29),
    .A2(net64),
    .B1(net34),
    .B2(net28),
    .X(_05460_));
 sky130_fd_sc_hd__and2b_1 _06329_ (.A_N(_05459_),
    .B(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__nand2_1 _06330_ (.A(net27),
    .B(net35),
    .Y(_05462_));
 sky130_fd_sc_hd__xnor2_1 _06331_ (.A(_05461_),
    .B(_05462_),
    .Y(_05463_));
 sky130_fd_sc_hd__o21ba_1 _06332_ (.A1(_05381_),
    .A2(_05383_),
    .B1_N(_05380_),
    .X(_05464_));
 sky130_fd_sc_hd__and2b_1 _06333_ (.A_N(_05464_),
    .B(_05463_),
    .X(_05465_));
 sky130_fd_sc_hd__xnor2_1 _06334_ (.A(_05463_),
    .B(_05464_),
    .Y(_05466_));
 sky130_fd_sc_hd__and2_1 _06335_ (.A(_05458_),
    .B(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__xnor2_1 _06336_ (.A(_05458_),
    .B(_05466_),
    .Y(_05468_));
 sky130_fd_sc_hd__a21o_1 _06337_ (.A1(_05401_),
    .A2(_05403_),
    .B1(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__nand3_1 _06338_ (.A(_05401_),
    .B(_05403_),
    .C(_05468_),
    .Y(_05470_));
 sky130_fd_sc_hd__o211ai_2 _06339_ (.A1(_05386_),
    .A2(_05388_),
    .B1(_05469_),
    .C1(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__a211o_1 _06340_ (.A1(_05469_),
    .A2(_05470_),
    .B1(_05386_),
    .C1(_05388_),
    .X(_05472_));
 sky130_fd_sc_hd__a31o_1 _06341_ (.A1(net29),
    .A2(net63),
    .A3(_05398_),
    .B1(_05396_),
    .X(_05473_));
 sky130_fd_sc_hd__o21bai_1 _06342_ (.A1(_05406_),
    .A2(_05408_),
    .B1_N(_05405_),
    .Y(_05474_));
 sky130_fd_sc_hd__nand4_1 _06343_ (.A(net61),
    .B(net62),
    .C(net31),
    .D(net32),
    .Y(_05475_));
 sky130_fd_sc_hd__a22o_1 _06344_ (.A1(net62),
    .A2(net31),
    .B1(net32),
    .B2(net61),
    .X(_05476_));
 sky130_fd_sc_hd__a22o_1 _06345_ (.A1(net30),
    .A2(net63),
    .B1(_05475_),
    .B2(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__nand4_1 _06346_ (.A(net30),
    .B(net63),
    .C(_05475_),
    .D(_05476_),
    .Y(_05478_));
 sky130_fd_sc_hd__and3_1 _06347_ (.A(_05474_),
    .B(_05477_),
    .C(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__a21o_1 _06348_ (.A1(_05477_),
    .A2(_05478_),
    .B1(_05474_),
    .X(_05480_));
 sky130_fd_sc_hd__and2b_1 _06349_ (.A_N(_05479_),
    .B(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__xor2_1 _06350_ (.A(_05473_),
    .B(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__and4_1 _06351_ (.A(net58),
    .B(net59),
    .C(net3),
    .D(net4),
    .X(_05483_));
 sky130_fd_sc_hd__a22oi_1 _06352_ (.A1(net59),
    .A2(net3),
    .B1(net4),
    .B2(net58),
    .Y(_05484_));
 sky130_fd_sc_hd__nor2_1 _06353_ (.A(_05483_),
    .B(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__nand2_1 _06354_ (.A(net60),
    .B(net2),
    .Y(_05486_));
 sky130_fd_sc_hd__xnor2_1 _06355_ (.A(_05485_),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__nand2_1 _06356_ (.A(net55),
    .B(net5),
    .Y(_05488_));
 sky130_fd_sc_hd__and4_1 _06357_ (.A(net33),
    .B(net44),
    .C(net6),
    .D(net7),
    .X(_05489_));
 sky130_fd_sc_hd__a22oi_2 _06358_ (.A1(net44),
    .A2(net6),
    .B1(net7),
    .B2(net33),
    .Y(_05490_));
 sky130_fd_sc_hd__or3_1 _06359_ (.A(_05488_),
    .B(_05489_),
    .C(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__o21ai_1 _06360_ (.A1(_05489_),
    .A2(_05490_),
    .B1(_05488_),
    .Y(_05492_));
 sky130_fd_sc_hd__o21bai_1 _06361_ (.A1(_05410_),
    .A2(_05412_),
    .B1_N(_05411_),
    .Y(_05493_));
 sky130_fd_sc_hd__nand3_1 _06362_ (.A(_05491_),
    .B(_05492_),
    .C(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__a21o_1 _06363_ (.A1(_05491_),
    .A2(_05492_),
    .B1(_05493_),
    .X(_05495_));
 sky130_fd_sc_hd__nand3_1 _06364_ (.A(_05487_),
    .B(_05494_),
    .C(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__a21o_1 _06365_ (.A1(_05494_),
    .A2(_05495_),
    .B1(_05487_),
    .X(_05497_));
 sky130_fd_sc_hd__a21bo_1 _06366_ (.A1(_05409_),
    .A2(_05417_),
    .B1_N(_05416_),
    .X(_05498_));
 sky130_fd_sc_hd__nand3_2 _06367_ (.A(_05496_),
    .B(_05497_),
    .C(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__a21o_1 _06368_ (.A1(_05496_),
    .A2(_05497_),
    .B1(_05498_),
    .X(_05500_));
 sky130_fd_sc_hd__and3_1 _06369_ (.A(_05482_),
    .B(_05499_),
    .C(_05500_),
    .X(_05501_));
 sky130_fd_sc_hd__nand3_1 _06370_ (.A(_05482_),
    .B(_05499_),
    .C(_05500_),
    .Y(_05502_));
 sky130_fd_sc_hd__a21oi_1 _06371_ (.A1(_05499_),
    .A2(_05500_),
    .B1(_05482_),
    .Y(_05503_));
 sky130_fd_sc_hd__a211o_1 _06372_ (.A1(_05421_),
    .A2(_05424_),
    .B1(_05501_),
    .C1(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__o211ai_2 _06373_ (.A1(_05501_),
    .A2(_05503_),
    .B1(_05421_),
    .C1(_05424_),
    .Y(_05505_));
 sky130_fd_sc_hd__and4_1 _06374_ (.A(_05471_),
    .B(_05472_),
    .C(_05504_),
    .D(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__nand4_1 _06375_ (.A(_05471_),
    .B(_05472_),
    .C(_05504_),
    .D(_05505_),
    .Y(_05507_));
 sky130_fd_sc_hd__a22oi_1 _06376_ (.A1(_05471_),
    .A2(_05472_),
    .B1(_05504_),
    .B2(_05505_),
    .Y(_05508_));
 sky130_fd_sc_hd__a211o_1 _06377_ (.A1(_05426_),
    .A2(_05429_),
    .B1(_05506_),
    .C1(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__inv_2 _06378_ (.A(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__o211ai_1 _06379_ (.A1(_05506_),
    .A2(_05508_),
    .B1(_05426_),
    .C1(_05429_),
    .Y(_05511_));
 sky130_fd_sc_hd__and3_1 _06380_ (.A(_05452_),
    .B(_05509_),
    .C(_05511_),
    .X(_05512_));
 sky130_fd_sc_hd__a21oi_1 _06381_ (.A1(_05509_),
    .A2(_05511_),
    .B1(_05452_),
    .Y(_05513_));
 sky130_fd_sc_hd__or2_1 _06382_ (.A(_05512_),
    .B(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__nand2_1 _06383_ (.A(_05431_),
    .B(_05433_),
    .Y(_05515_));
 sky130_fd_sc_hd__a211oi_1 _06384_ (.A1(_05431_),
    .A2(_05433_),
    .B1(_05512_),
    .C1(_05513_),
    .Y(_05516_));
 sky130_fd_sc_hd__xnor2_1 _06385_ (.A(_05514_),
    .B(_05515_),
    .Y(_05517_));
 sky130_fd_sc_hd__a211oi_1 _06386_ (.A1(_05431_),
    .A2(_05514_),
    .B1(_05516_),
    .C1(_05371_),
    .Y(_05518_));
 sky130_fd_sc_hd__xnor2_1 _06387_ (.A(_05371_),
    .B(_05517_),
    .Y(_05519_));
 sky130_fd_sc_hd__and2_1 _06388_ (.A(_05437_),
    .B(_05519_),
    .X(_05520_));
 sky130_fd_sc_hd__xor2_2 _06389_ (.A(_05437_),
    .B(_05519_),
    .X(_05521_));
 sky130_fd_sc_hd__o21a_1 _06390_ (.A1(_05365_),
    .A2(_05441_),
    .B1(_05439_),
    .X(_05522_));
 sky130_fd_sc_hd__xnor2_1 _06391_ (.A(_05521_),
    .B(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__xor2_1 _06392_ (.A(_05445_),
    .B(_05523_),
    .X(net71));
 sky130_fd_sc_hd__a22o_2 _06393_ (.A1(_05442_),
    .A2(_05521_),
    .B1(_05523_),
    .B2(_05445_),
    .X(_05524_));
 sky130_fd_sc_hd__nand2b_1 _06394_ (.A_N(_05439_),
    .B(_05521_),
    .Y(_05525_));
 sky130_fd_sc_hd__and4_1 _06395_ (.A(net12),
    .B(net1),
    .C(net39),
    .D(net40),
    .X(_05526_));
 sky130_fd_sc_hd__nand4_1 _06396_ (.A(net12),
    .B(net1),
    .C(net39),
    .D(net40),
    .Y(_05527_));
 sky130_fd_sc_hd__a22o_1 _06397_ (.A1(net12),
    .A2(net39),
    .B1(net40),
    .B2(net1),
    .X(_05528_));
 sky130_fd_sc_hd__o211a_1 _06398_ (.A1(_05453_),
    .A2(_05457_),
    .B1(_05527_),
    .C1(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__a211oi_1 _06399_ (.A1(_05527_),
    .A2(_05528_),
    .B1(_05453_),
    .C1(_05457_),
    .Y(_05530_));
 sky130_fd_sc_hd__nor2_1 _06400_ (.A(_05529_),
    .B(_05530_),
    .Y(_05531_));
 sky130_fd_sc_hd__nand2_1 _06401_ (.A(_05448_),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__or2_1 _06402_ (.A(_05448_),
    .B(_05531_),
    .X(_05533_));
 sky130_fd_sc_hd__nand2_1 _06403_ (.A(_05532_),
    .B(_05533_),
    .Y(_05534_));
 sky130_fd_sc_hd__a21oi_1 _06404_ (.A1(_05469_),
    .A2(_05471_),
    .B1(_05534_),
    .Y(_05535_));
 sky130_fd_sc_hd__and3_1 _06405_ (.A(_05469_),
    .B(_05471_),
    .C(_05534_),
    .X(_05536_));
 sky130_fd_sc_hd__nor2_1 _06406_ (.A(_05535_),
    .B(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__a21o_1 _06407_ (.A1(_05473_),
    .A2(_05480_),
    .B1(_05479_),
    .X(_05538_));
 sky130_fd_sc_hd__and4_1 _06408_ (.A(net27),
    .B(net26),
    .C(net36),
    .D(net37),
    .X(_05539_));
 sky130_fd_sc_hd__a22o_1 _06409_ (.A1(net27),
    .A2(net36),
    .B1(net37),
    .B2(net26),
    .X(_05540_));
 sky130_fd_sc_hd__and2b_1 _06410_ (.A_N(_05539_),
    .B(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__nand2_1 _06411_ (.A(net23),
    .B(net38),
    .Y(_05542_));
 sky130_fd_sc_hd__xnor2_1 _06412_ (.A(_05541_),
    .B(_05542_),
    .Y(_05543_));
 sky130_fd_sc_hd__nand4_1 _06413_ (.A(net29),
    .B(net30),
    .C(net64),
    .D(net34),
    .Y(_05544_));
 sky130_fd_sc_hd__a22o_1 _06414_ (.A1(net30),
    .A2(net64),
    .B1(net34),
    .B2(net29),
    .X(_05545_));
 sky130_fd_sc_hd__and2_1 _06415_ (.A(net28),
    .B(net35),
    .X(_05546_));
 sky130_fd_sc_hd__a21o_1 _06416_ (.A1(_05544_),
    .A2(_05545_),
    .B1(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__nand3_1 _06417_ (.A(_05544_),
    .B(_05545_),
    .C(_05546_),
    .Y(_05548_));
 sky130_fd_sc_hd__a31o_1 _06418_ (.A1(net27),
    .A2(net35),
    .A3(_05460_),
    .B1(_05459_),
    .X(_05549_));
 sky130_fd_sc_hd__nand3_1 _06419_ (.A(_05547_),
    .B(_05548_),
    .C(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__a21o_1 _06420_ (.A1(_05547_),
    .A2(_05548_),
    .B1(_05549_),
    .X(_05551_));
 sky130_fd_sc_hd__nand3_1 _06421_ (.A(_05543_),
    .B(_05550_),
    .C(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__a21o_1 _06422_ (.A1(_05550_),
    .A2(_05551_),
    .B1(_05543_),
    .X(_05553_));
 sky130_fd_sc_hd__nand3_2 _06423_ (.A(_05538_),
    .B(_05552_),
    .C(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__a21o_1 _06424_ (.A1(_05552_),
    .A2(_05553_),
    .B1(_05538_),
    .X(_05555_));
 sky130_fd_sc_hd__o211ai_2 _06425_ (.A1(_05465_),
    .A2(_05467_),
    .B1(_05554_),
    .C1(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__a211o_1 _06426_ (.A1(_05554_),
    .A2(_05555_),
    .B1(_05465_),
    .C1(_05467_),
    .X(_05557_));
 sky130_fd_sc_hd__nand2_1 _06427_ (.A(_05556_),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__nand2_1 _06428_ (.A(_05475_),
    .B(_05478_),
    .Y(_05559_));
 sky130_fd_sc_hd__o21bai_1 _06429_ (.A1(_05484_),
    .A2(_05486_),
    .B1_N(_05483_),
    .Y(_05560_));
 sky130_fd_sc_hd__nand4_1 _06430_ (.A(net61),
    .B(net62),
    .C(net2),
    .D(net32),
    .Y(_05561_));
 sky130_fd_sc_hd__a22o_1 _06431_ (.A1(net61),
    .A2(net2),
    .B1(net32),
    .B2(net62),
    .X(_05562_));
 sky130_fd_sc_hd__a22o_1 _06432_ (.A1(net31),
    .A2(net63),
    .B1(_05561_),
    .B2(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__nand4_1 _06433_ (.A(net31),
    .B(net63),
    .C(_05561_),
    .D(_05562_),
    .Y(_05564_));
 sky130_fd_sc_hd__and3_1 _06434_ (.A(_05560_),
    .B(_05563_),
    .C(_05564_),
    .X(_05565_));
 sky130_fd_sc_hd__a21o_1 _06435_ (.A1(_05563_),
    .A2(_05564_),
    .B1(_05560_),
    .X(_05566_));
 sky130_fd_sc_hd__and2b_1 _06436_ (.A_N(_05565_),
    .B(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__xor2_1 _06437_ (.A(_05559_),
    .B(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__and4_1 _06438_ (.A(net58),
    .B(net59),
    .C(net4),
    .D(net5),
    .X(_05569_));
 sky130_fd_sc_hd__a22oi_1 _06439_ (.A1(net59),
    .A2(net4),
    .B1(net5),
    .B2(net58),
    .Y(_05570_));
 sky130_fd_sc_hd__nor2_1 _06440_ (.A(_05569_),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__nand2_1 _06441_ (.A(net60),
    .B(net3),
    .Y(_05572_));
 sky130_fd_sc_hd__xnor2_1 _06442_ (.A(_05571_),
    .B(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__nand2_1 _06443_ (.A(net55),
    .B(net6),
    .Y(_05574_));
 sky130_fd_sc_hd__and4_1 _06444_ (.A(net33),
    .B(net44),
    .C(net7),
    .D(net8),
    .X(_05575_));
 sky130_fd_sc_hd__a22oi_2 _06445_ (.A1(net44),
    .A2(net7),
    .B1(net8),
    .B2(net33),
    .Y(_05576_));
 sky130_fd_sc_hd__or3_1 _06446_ (.A(_05574_),
    .B(_05575_),
    .C(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__o21ai_1 _06447_ (.A1(_05575_),
    .A2(_05576_),
    .B1(_05574_),
    .Y(_05578_));
 sky130_fd_sc_hd__o21bai_1 _06448_ (.A1(_05488_),
    .A2(_05490_),
    .B1_N(_05489_),
    .Y(_05579_));
 sky130_fd_sc_hd__nand3_1 _06449_ (.A(_05577_),
    .B(_05578_),
    .C(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__a21o_1 _06450_ (.A1(_05577_),
    .A2(_05578_),
    .B1(_05579_),
    .X(_05581_));
 sky130_fd_sc_hd__nand3_1 _06451_ (.A(_05573_),
    .B(_05580_),
    .C(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__a21o_1 _06452_ (.A1(_05580_),
    .A2(_05581_),
    .B1(_05573_),
    .X(_05583_));
 sky130_fd_sc_hd__a21bo_1 _06453_ (.A1(_05487_),
    .A2(_05495_),
    .B1_N(_05494_),
    .X(_05584_));
 sky130_fd_sc_hd__nand3_2 _06454_ (.A(_05582_),
    .B(_05583_),
    .C(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__a21o_1 _06455_ (.A1(_05582_),
    .A2(_05583_),
    .B1(_05584_),
    .X(_05586_));
 sky130_fd_sc_hd__and3_1 _06456_ (.A(_05568_),
    .B(_05585_),
    .C(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__nand3_1 _06457_ (.A(_05568_),
    .B(_05585_),
    .C(_05586_),
    .Y(_05588_));
 sky130_fd_sc_hd__a21oi_1 _06458_ (.A1(_05585_),
    .A2(_05586_),
    .B1(_05568_),
    .Y(_05589_));
 sky130_fd_sc_hd__a211oi_2 _06459_ (.A1(_05499_),
    .A2(_05502_),
    .B1(_05587_),
    .C1(_05589_),
    .Y(_05590_));
 sky130_fd_sc_hd__o211a_1 _06460_ (.A1(_05587_),
    .A2(_05589_),
    .B1(_05499_),
    .C1(_05502_),
    .X(_05591_));
 sky130_fd_sc_hd__nor3_2 _06461_ (.A(_05558_),
    .B(_05590_),
    .C(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__o21a_1 _06462_ (.A1(_05590_),
    .A2(_05591_),
    .B1(_05558_),
    .X(_05593_));
 sky130_fd_sc_hd__a211o_1 _06463_ (.A1(_05504_),
    .A2(_05507_),
    .B1(_05592_),
    .C1(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__o211ai_2 _06464_ (.A1(_05592_),
    .A2(_05593_),
    .B1(_05504_),
    .C1(_05507_),
    .Y(_05595_));
 sky130_fd_sc_hd__nand3_2 _06465_ (.A(_05537_),
    .B(_05594_),
    .C(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__a21o_1 _06466_ (.A1(_05594_),
    .A2(_05595_),
    .B1(_05537_),
    .X(_05597_));
 sky130_fd_sc_hd__o211ai_4 _06467_ (.A1(_05510_),
    .A2(_05512_),
    .B1(_05596_),
    .C1(_05597_),
    .Y(_05598_));
 sky130_fd_sc_hd__a211o_1 _06468_ (.A1(_05596_),
    .A2(_05597_),
    .B1(_05510_),
    .C1(_05512_),
    .X(_05599_));
 sky130_fd_sc_hd__nand3_2 _06469_ (.A(_05450_),
    .B(_05598_),
    .C(_05599_),
    .Y(_05600_));
 sky130_fd_sc_hd__a21o_1 _06470_ (.A1(_05598_),
    .A2(_05599_),
    .B1(_05450_),
    .X(_05601_));
 sky130_fd_sc_hd__o211a_1 _06471_ (.A1(_05516_),
    .A2(_05518_),
    .B1(_05600_),
    .C1(_05601_),
    .X(_05602_));
 sky130_fd_sc_hd__a211oi_1 _06472_ (.A1(_05600_),
    .A2(_05601_),
    .B1(_05516_),
    .C1(_05518_),
    .Y(_05603_));
 sky130_fd_sc_hd__nor2_1 _06473_ (.A(_05602_),
    .B(_05603_),
    .Y(_05604_));
 sky130_fd_sc_hd__inv_2 _06474_ (.A(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__nand3b_1 _06475_ (.A_N(_05520_),
    .B(_05525_),
    .C(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__nand2_1 _06476_ (.A(_05520_),
    .B(_05604_),
    .Y(_05607_));
 sky130_fd_sc_hd__o211a_1 _06477_ (.A1(_05525_),
    .A2(_05605_),
    .B1(_05606_),
    .C1(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__xor2_1 _06478_ (.A(_05524_),
    .B(_05608_),
    .X(net72));
 sky130_fd_sc_hd__o2bb2a_1 _06479_ (.A1_N(_05524_),
    .A2_N(_05608_),
    .B1(_05605_),
    .B2(_05525_),
    .X(_05609_));
 sky130_fd_sc_hd__a31o_1 _06480_ (.A1(net23),
    .A2(net38),
    .A3(_05540_),
    .B1(_05539_),
    .X(_05610_));
 sky130_fd_sc_hd__and4_1 _06481_ (.A(net23),
    .B(net12),
    .C(net39),
    .D(net40),
    .X(_05611_));
 sky130_fd_sc_hd__a22oi_1 _06482_ (.A1(net23),
    .A2(net39),
    .B1(net40),
    .B2(net12),
    .Y(_05612_));
 sky130_fd_sc_hd__and4bb_1 _06483_ (.A_N(_05611_),
    .B_N(_05612_),
    .C(net1),
    .D(net41),
    .X(_05613_));
 sky130_fd_sc_hd__o2bb2a_1 _06484_ (.A1_N(net1),
    .A2_N(net41),
    .B1(_05611_),
    .B2(_05612_),
    .X(_05614_));
 sky130_fd_sc_hd__nor2_1 _06485_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__or2_1 _06486_ (.A(_05610_),
    .B(_05615_),
    .X(_05616_));
 sky130_fd_sc_hd__and2_1 _06487_ (.A(_05610_),
    .B(_05615_),
    .X(_05617_));
 sky130_fd_sc_hd__nand2_1 _06488_ (.A(_05610_),
    .B(_05615_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand2_1 _06489_ (.A(_05616_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__nor2_1 _06490_ (.A(_05526_),
    .B(_05529_),
    .Y(_05620_));
 sky130_fd_sc_hd__xnor2_1 _06491_ (.A(_05619_),
    .B(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__and3_1 _06492_ (.A(_05554_),
    .B(_05556_),
    .C(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__a21o_1 _06493_ (.A1(_05554_),
    .A2(_05556_),
    .B1(_05621_),
    .X(_05623_));
 sky130_fd_sc_hd__nand2b_1 _06494_ (.A_N(_05622_),
    .B(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__xor2_1 _06495_ (.A(_05532_),
    .B(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__nand2_1 _06496_ (.A(_05550_),
    .B(_05552_),
    .Y(_05626_));
 sky130_fd_sc_hd__a21o_1 _06497_ (.A1(_05559_),
    .A2(_05566_),
    .B1(_05565_),
    .X(_05627_));
 sky130_fd_sc_hd__nand2_1 _06498_ (.A(net26),
    .B(net38),
    .Y(_05628_));
 sky130_fd_sc_hd__and4_1 _06499_ (.A(net28),
    .B(net27),
    .C(net36),
    .D(net37),
    .X(_05629_));
 sky130_fd_sc_hd__a22oi_1 _06500_ (.A1(net28),
    .A2(net36),
    .B1(net37),
    .B2(net27),
    .Y(_05630_));
 sky130_fd_sc_hd__nor2_1 _06501_ (.A(_05629_),
    .B(_05630_),
    .Y(_05631_));
 sky130_fd_sc_hd__xnor2_1 _06502_ (.A(_05628_),
    .B(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__nand2_1 _06503_ (.A(net29),
    .B(net35),
    .Y(_05633_));
 sky130_fd_sc_hd__nand4_1 _06504_ (.A(net30),
    .B(net31),
    .C(net64),
    .D(net34),
    .Y(_05634_));
 sky130_fd_sc_hd__a22o_1 _06505_ (.A1(net31),
    .A2(net64),
    .B1(net34),
    .B2(net30),
    .X(_05635_));
 sky130_fd_sc_hd__nand3b_1 _06506_ (.A_N(_05633_),
    .B(_05634_),
    .C(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hd__a21bo_1 _06507_ (.A1(_05634_),
    .A2(_05635_),
    .B1_N(_05633_),
    .X(_05637_));
 sky130_fd_sc_hd__a21bo_1 _06508_ (.A1(_05545_),
    .A2(_05546_),
    .B1_N(_05544_),
    .X(_05638_));
 sky130_fd_sc_hd__nand3_1 _06509_ (.A(_05636_),
    .B(_05637_),
    .C(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__a21o_1 _06510_ (.A1(_05636_),
    .A2(_05637_),
    .B1(_05638_),
    .X(_05640_));
 sky130_fd_sc_hd__nand3_1 _06511_ (.A(_05632_),
    .B(_05639_),
    .C(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__a21o_1 _06512_ (.A1(_05639_),
    .A2(_05640_),
    .B1(_05632_),
    .X(_05642_));
 sky130_fd_sc_hd__nand3_1 _06513_ (.A(_05627_),
    .B(_05641_),
    .C(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__a21o_1 _06514_ (.A1(_05641_),
    .A2(_05642_),
    .B1(_05627_),
    .X(_05644_));
 sky130_fd_sc_hd__and3_1 _06515_ (.A(_05626_),
    .B(_05643_),
    .C(_05644_),
    .X(_05645_));
 sky130_fd_sc_hd__a21oi_1 _06516_ (.A1(_05643_),
    .A2(_05644_),
    .B1(_05626_),
    .Y(_05646_));
 sky130_fd_sc_hd__or2_1 _06517_ (.A(_05645_),
    .B(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__nand2_1 _06518_ (.A(_05561_),
    .B(_05564_),
    .Y(_05648_));
 sky130_fd_sc_hd__o21ba_1 _06519_ (.A1(_05570_),
    .A2(_05572_),
    .B1_N(_05569_),
    .X(_05649_));
 sky130_fd_sc_hd__nand2_1 _06520_ (.A(net63),
    .B(net32),
    .Y(_05650_));
 sky130_fd_sc_hd__and4_1 _06521_ (.A(net61),
    .B(net62),
    .C(net2),
    .D(net3),
    .X(_05651_));
 sky130_fd_sc_hd__a22oi_1 _06522_ (.A1(net62),
    .A2(net2),
    .B1(net3),
    .B2(net61),
    .Y(_05652_));
 sky130_fd_sc_hd__nor2_1 _06523_ (.A(_05651_),
    .B(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__xnor2_1 _06524_ (.A(_05650_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand2b_1 _06525_ (.A_N(_05649_),
    .B(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__xnor2_1 _06526_ (.A(_05649_),
    .B(_05654_),
    .Y(_05656_));
 sky130_fd_sc_hd__nand2_1 _06527_ (.A(_05648_),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__xor2_1 _06528_ (.A(_05648_),
    .B(_05656_),
    .X(_05658_));
 sky130_fd_sc_hd__nand2_1 _06529_ (.A(net60),
    .B(net4),
    .Y(_05659_));
 sky130_fd_sc_hd__and4_1 _06530_ (.A(net58),
    .B(net59),
    .C(net5),
    .D(net6),
    .X(_05660_));
 sky130_fd_sc_hd__a22oi_1 _06531_ (.A1(net59),
    .A2(net5),
    .B1(net6),
    .B2(net58),
    .Y(_05661_));
 sky130_fd_sc_hd__nor2_1 _06532_ (.A(_05660_),
    .B(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__xnor2_1 _06533_ (.A(_05659_),
    .B(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__nand2_1 _06534_ (.A(net55),
    .B(net7),
    .Y(_05664_));
 sky130_fd_sc_hd__and4_1 _06535_ (.A(net33),
    .B(net44),
    .C(net8),
    .D(net9),
    .X(_05665_));
 sky130_fd_sc_hd__a22oi_2 _06536_ (.A1(net44),
    .A2(net8),
    .B1(net9),
    .B2(net33),
    .Y(_05666_));
 sky130_fd_sc_hd__or3_1 _06537_ (.A(_05664_),
    .B(_05665_),
    .C(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__o21ai_1 _06538_ (.A1(_05665_),
    .A2(_05666_),
    .B1(_05664_),
    .Y(_05668_));
 sky130_fd_sc_hd__o21bai_1 _06539_ (.A1(_05574_),
    .A2(_05576_),
    .B1_N(_05575_),
    .Y(_05669_));
 sky130_fd_sc_hd__nand3_1 _06540_ (.A(_05667_),
    .B(_05668_),
    .C(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__a21o_1 _06541_ (.A1(_05667_),
    .A2(_05668_),
    .B1(_05669_),
    .X(_05671_));
 sky130_fd_sc_hd__nand3_1 _06542_ (.A(_05663_),
    .B(_05670_),
    .C(_05671_),
    .Y(_05672_));
 sky130_fd_sc_hd__a21o_1 _06543_ (.A1(_05670_),
    .A2(_05671_),
    .B1(_05663_),
    .X(_05673_));
 sky130_fd_sc_hd__a21bo_1 _06544_ (.A1(_05573_),
    .A2(_05581_),
    .B1_N(_05580_),
    .X(_05674_));
 sky130_fd_sc_hd__nand3_2 _06545_ (.A(_05672_),
    .B(_05673_),
    .C(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__a21o_1 _06546_ (.A1(_05672_),
    .A2(_05673_),
    .B1(_05674_),
    .X(_05676_));
 sky130_fd_sc_hd__and3_1 _06547_ (.A(_05658_),
    .B(_05675_),
    .C(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__nand3_1 _06548_ (.A(_05658_),
    .B(_05675_),
    .C(_05676_),
    .Y(_05678_));
 sky130_fd_sc_hd__a21oi_1 _06549_ (.A1(_05675_),
    .A2(_05676_),
    .B1(_05658_),
    .Y(_05679_));
 sky130_fd_sc_hd__a211oi_2 _06550_ (.A1(_05585_),
    .A2(_05588_),
    .B1(_05677_),
    .C1(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__o211a_1 _06551_ (.A1(_05677_),
    .A2(_05679_),
    .B1(_05585_),
    .C1(_05588_),
    .X(_05681_));
 sky130_fd_sc_hd__nor3_1 _06552_ (.A(_05647_),
    .B(_05680_),
    .C(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__or3_1 _06553_ (.A(_05647_),
    .B(_05680_),
    .C(_05681_),
    .X(_05683_));
 sky130_fd_sc_hd__o21ai_1 _06554_ (.A1(_05680_),
    .A2(_05681_),
    .B1(_05647_),
    .Y(_05684_));
 sky130_fd_sc_hd__o211ai_2 _06555_ (.A1(_05590_),
    .A2(_05592_),
    .B1(_05683_),
    .C1(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__a211o_1 _06556_ (.A1(_05683_),
    .A2(_05684_),
    .B1(_05590_),
    .C1(_05592_),
    .X(_05686_));
 sky130_fd_sc_hd__and3_1 _06557_ (.A(_05625_),
    .B(_05685_),
    .C(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__a21oi_1 _06558_ (.A1(_05685_),
    .A2(_05686_),
    .B1(_05625_),
    .Y(_05688_));
 sky130_fd_sc_hd__a211o_1 _06559_ (.A1(_05594_),
    .A2(_05596_),
    .B1(_05687_),
    .C1(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__inv_2 _06560_ (.A(_05689_),
    .Y(_05690_));
 sky130_fd_sc_hd__o211ai_1 _06561_ (.A1(_05687_),
    .A2(_05688_),
    .B1(_05594_),
    .C1(_05596_),
    .Y(_05691_));
 sky130_fd_sc_hd__and3_1 _06562_ (.A(_05535_),
    .B(_05689_),
    .C(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__a21oi_1 _06563_ (.A1(_05689_),
    .A2(_05691_),
    .B1(_05535_),
    .Y(_05693_));
 sky130_fd_sc_hd__a211o_1 _06564_ (.A1(_05598_),
    .A2(_05600_),
    .B1(_05692_),
    .C1(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__o211ai_1 _06565_ (.A1(_05692_),
    .A2(_05693_),
    .B1(_05598_),
    .C1(_05600_),
    .Y(_05695_));
 sky130_fd_sc_hd__and3_1 _06566_ (.A(_05602_),
    .B(_05694_),
    .C(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__a21oi_1 _06567_ (.A1(_05694_),
    .A2(_05695_),
    .B1(_05602_),
    .Y(_05697_));
 sky130_fd_sc_hd__nor2_1 _06568_ (.A(_05696_),
    .B(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__or3_1 _06569_ (.A(_05607_),
    .B(_05696_),
    .C(_05697_),
    .X(_05699_));
 sky130_fd_sc_hd__xnor2_1 _06570_ (.A(_05607_),
    .B(_05698_),
    .Y(_05700_));
 sky130_fd_sc_hd__xnor2_1 _06571_ (.A(_05609_),
    .B(_05700_),
    .Y(net73));
 sky130_fd_sc_hd__nor2_1 _06572_ (.A(_05690_),
    .B(_05692_),
    .Y(_05701_));
 sky130_fd_sc_hd__o21a_1 _06573_ (.A1(_05532_),
    .A2(_05622_),
    .B1(_05623_),
    .X(_05702_));
 sky130_fd_sc_hd__and3b_1 _06574_ (.A_N(_05617_),
    .B(_05529_),
    .C(_05616_),
    .X(_05703_));
 sky130_fd_sc_hd__a31o_1 _06575_ (.A1(_05627_),
    .A2(_05641_),
    .A3(_05642_),
    .B1(_05645_),
    .X(_05704_));
 sky130_fd_sc_hd__or2_1 _06576_ (.A(_05611_),
    .B(_05613_),
    .X(_05705_));
 sky130_fd_sc_hd__o21ba_1 _06577_ (.A1(_05628_),
    .A2(_05630_),
    .B1_N(_05629_),
    .X(_05706_));
 sky130_fd_sc_hd__and4_1 _06578_ (.A(net26),
    .B(net23),
    .C(net39),
    .D(net40),
    .X(_05707_));
 sky130_fd_sc_hd__a22oi_1 _06579_ (.A1(net26),
    .A2(net39),
    .B1(net40),
    .B2(net23),
    .Y(_05708_));
 sky130_fd_sc_hd__nor2_1 _06580_ (.A(_05707_),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__nand2_1 _06581_ (.A(net12),
    .B(net41),
    .Y(_05710_));
 sky130_fd_sc_hd__xnor2_1 _06582_ (.A(_05709_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__nand2b_1 _06583_ (.A_N(_05706_),
    .B(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__xnor2_1 _06584_ (.A(_05706_),
    .B(_05711_),
    .Y(_05713_));
 sky130_fd_sc_hd__nand2_1 _06585_ (.A(_05705_),
    .B(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__xnor2_1 _06586_ (.A(_05705_),
    .B(_05713_),
    .Y(_05715_));
 sky130_fd_sc_hd__o21ai_1 _06587_ (.A1(_05526_),
    .A2(_05617_),
    .B1(_05616_),
    .Y(_05716_));
 sky130_fd_sc_hd__xor2_1 _06588_ (.A(_05715_),
    .B(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__nand2_1 _06589_ (.A(net1),
    .B(net42),
    .Y(_05718_));
 sky130_fd_sc_hd__and3_1 _06590_ (.A(net1),
    .B(net42),
    .C(_05717_),
    .X(_05719_));
 sky130_fd_sc_hd__xor2_1 _06591_ (.A(_05717_),
    .B(_05718_),
    .X(_05720_));
 sky130_fd_sc_hd__and2b_1 _06592_ (.A_N(_05720_),
    .B(_05704_),
    .X(_05721_));
 sky130_fd_sc_hd__xnor2_1 _06593_ (.A(_05704_),
    .B(_05720_),
    .Y(_05722_));
 sky130_fd_sc_hd__xnor2_1 _06594_ (.A(_05703_),
    .B(_05722_),
    .Y(_05723_));
 sky130_fd_sc_hd__nand2_1 _06595_ (.A(_05639_),
    .B(_05641_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand2_1 _06596_ (.A(net27),
    .B(net38),
    .Y(_05725_));
 sky130_fd_sc_hd__and4_1 _06597_ (.A(net28),
    .B(net29),
    .C(net36),
    .D(net37),
    .X(_05726_));
 sky130_fd_sc_hd__a22oi_1 _06598_ (.A1(net29),
    .A2(net36),
    .B1(net37),
    .B2(net28),
    .Y(_05727_));
 sky130_fd_sc_hd__nor2_1 _06599_ (.A(_05726_),
    .B(_05727_),
    .Y(_05728_));
 sky130_fd_sc_hd__xnor2_1 _06600_ (.A(_05725_),
    .B(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__nand2_1 _06601_ (.A(net30),
    .B(net35),
    .Y(_05730_));
 sky130_fd_sc_hd__and4_1 _06602_ (.A(net31),
    .B(net32),
    .C(net64),
    .D(net34),
    .X(_05731_));
 sky130_fd_sc_hd__a22oi_1 _06603_ (.A1(net32),
    .A2(net64),
    .B1(net34),
    .B2(net31),
    .Y(_05732_));
 sky130_fd_sc_hd__nor2_1 _06604_ (.A(_05731_),
    .B(_05732_),
    .Y(_05733_));
 sky130_fd_sc_hd__xnor2_1 _06605_ (.A(_05730_),
    .B(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__nand2_1 _06606_ (.A(_05634_),
    .B(_05636_),
    .Y(_05735_));
 sky130_fd_sc_hd__and2_1 _06607_ (.A(_05734_),
    .B(_05735_),
    .X(_05736_));
 sky130_fd_sc_hd__xor2_1 _06608_ (.A(_05734_),
    .B(_05735_),
    .X(_05737_));
 sky130_fd_sc_hd__and2_1 _06609_ (.A(_05729_),
    .B(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__xnor2_1 _06610_ (.A(_05729_),
    .B(_05737_),
    .Y(_05739_));
 sky130_fd_sc_hd__a21o_1 _06611_ (.A1(_05655_),
    .A2(_05657_),
    .B1(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__nand3_1 _06612_ (.A(_05655_),
    .B(_05657_),
    .C(_05739_),
    .Y(_05741_));
 sky130_fd_sc_hd__and3_1 _06613_ (.A(_05724_),
    .B(_05740_),
    .C(_05741_),
    .X(_05742_));
 sky130_fd_sc_hd__nand3_1 _06614_ (.A(_05724_),
    .B(_05740_),
    .C(_05741_),
    .Y(_05743_));
 sky130_fd_sc_hd__a21oi_1 _06615_ (.A1(_05740_),
    .A2(_05741_),
    .B1(_05724_),
    .Y(_05744_));
 sky130_fd_sc_hd__o21ba_1 _06616_ (.A1(_05650_),
    .A2(_05652_),
    .B1_N(_05651_),
    .X(_05745_));
 sky130_fd_sc_hd__o21ba_1 _06617_ (.A1(_05659_),
    .A2(_05661_),
    .B1_N(_05660_),
    .X(_05746_));
 sky130_fd_sc_hd__nand2_1 _06618_ (.A(net63),
    .B(net2),
    .Y(_05747_));
 sky130_fd_sc_hd__and4_1 _06619_ (.A(net61),
    .B(net62),
    .C(net3),
    .D(net4),
    .X(_05748_));
 sky130_fd_sc_hd__a22oi_1 _06620_ (.A1(net62),
    .A2(net3),
    .B1(net4),
    .B2(net61),
    .Y(_05749_));
 sky130_fd_sc_hd__nor2_1 _06621_ (.A(_05748_),
    .B(_05749_),
    .Y(_05750_));
 sky130_fd_sc_hd__xnor2_1 _06622_ (.A(_05747_),
    .B(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__nand2b_1 _06623_ (.A_N(_05746_),
    .B(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__xnor2_1 _06624_ (.A(_05746_),
    .B(_05751_),
    .Y(_05753_));
 sky130_fd_sc_hd__nand2b_1 _06625_ (.A_N(_05745_),
    .B(_05753_),
    .Y(_00000_));
 sky130_fd_sc_hd__xnor2_1 _06626_ (.A(_05745_),
    .B(_05753_),
    .Y(_00001_));
 sky130_fd_sc_hd__nand2_1 _06627_ (.A(net60),
    .B(net5),
    .Y(_00002_));
 sky130_fd_sc_hd__and4_1 _06628_ (.A(net58),
    .B(net59),
    .C(net6),
    .D(net7),
    .X(_00003_));
 sky130_fd_sc_hd__a22oi_1 _06629_ (.A1(net59),
    .A2(net6),
    .B1(net7),
    .B2(net58),
    .Y(_00004_));
 sky130_fd_sc_hd__nor2_1 _06630_ (.A(_00003_),
    .B(_00004_),
    .Y(_00005_));
 sky130_fd_sc_hd__xnor2_1 _06631_ (.A(_00002_),
    .B(_00005_),
    .Y(_00006_));
 sky130_fd_sc_hd__nand2_1 _06632_ (.A(net55),
    .B(net8),
    .Y(_00007_));
 sky130_fd_sc_hd__and4_1 _06633_ (.A(net33),
    .B(net44),
    .C(net9),
    .D(net10),
    .X(_00008_));
 sky130_fd_sc_hd__a22oi_2 _06634_ (.A1(net44),
    .A2(net9),
    .B1(net10),
    .B2(net33),
    .Y(_00009_));
 sky130_fd_sc_hd__or3_1 _06635_ (.A(_00007_),
    .B(_00008_),
    .C(_00009_),
    .X(_00010_));
 sky130_fd_sc_hd__o21ai_1 _06636_ (.A1(_00008_),
    .A2(_00009_),
    .B1(_00007_),
    .Y(_00011_));
 sky130_fd_sc_hd__o21bai_1 _06637_ (.A1(_05664_),
    .A2(_05666_),
    .B1_N(_05665_),
    .Y(_00012_));
 sky130_fd_sc_hd__nand3_1 _06638_ (.A(_00010_),
    .B(_00011_),
    .C(_00012_),
    .Y(_00013_));
 sky130_fd_sc_hd__a21o_1 _06639_ (.A1(_00010_),
    .A2(_00011_),
    .B1(_00012_),
    .X(_00014_));
 sky130_fd_sc_hd__nand3_1 _06640_ (.A(_00006_),
    .B(_00013_),
    .C(_00014_),
    .Y(_00015_));
 sky130_fd_sc_hd__a21o_1 _06641_ (.A1(_00013_),
    .A2(_00014_),
    .B1(_00006_),
    .X(_00016_));
 sky130_fd_sc_hd__a21bo_1 _06642_ (.A1(_05663_),
    .A2(_05671_),
    .B1_N(_05670_),
    .X(_00017_));
 sky130_fd_sc_hd__nand3_4 _06643_ (.A(_00015_),
    .B(_00016_),
    .C(_00017_),
    .Y(_00018_));
 sky130_fd_sc_hd__a21o_1 _06644_ (.A1(_00015_),
    .A2(_00016_),
    .B1(_00017_),
    .X(_00019_));
 sky130_fd_sc_hd__and3_1 _06645_ (.A(_00001_),
    .B(_00018_),
    .C(_00019_),
    .X(_00020_));
 sky130_fd_sc_hd__nand3_2 _06646_ (.A(_00001_),
    .B(_00018_),
    .C(_00019_),
    .Y(_00021_));
 sky130_fd_sc_hd__a21oi_1 _06647_ (.A1(_00018_),
    .A2(_00019_),
    .B1(_00001_),
    .Y(_00022_));
 sky130_fd_sc_hd__a211oi_2 _06648_ (.A1(_05675_),
    .A2(_05678_),
    .B1(_00020_),
    .C1(_00022_),
    .Y(_00023_));
 sky130_fd_sc_hd__o211a_1 _06649_ (.A1(_00020_),
    .A2(_00022_),
    .B1(_05675_),
    .C1(_05678_),
    .X(_00024_));
 sky130_fd_sc_hd__nor4_1 _06650_ (.A(_05742_),
    .B(_05744_),
    .C(_00023_),
    .D(_00024_),
    .Y(_00025_));
 sky130_fd_sc_hd__or4_1 _06651_ (.A(_05742_),
    .B(_05744_),
    .C(_00023_),
    .D(_00024_),
    .X(_00026_));
 sky130_fd_sc_hd__o22ai_1 _06652_ (.A1(_05742_),
    .A2(_05744_),
    .B1(_00023_),
    .B2(_00024_),
    .Y(_00027_));
 sky130_fd_sc_hd__o211a_1 _06653_ (.A1(_05680_),
    .A2(_05682_),
    .B1(_00026_),
    .C1(_00027_),
    .X(_00028_));
 sky130_fd_sc_hd__a211oi_1 _06654_ (.A1(_00026_),
    .A2(_00027_),
    .B1(_05680_),
    .C1(_05682_),
    .Y(_00029_));
 sky130_fd_sc_hd__or3_1 _06655_ (.A(_05723_),
    .B(_00028_),
    .C(_00029_),
    .X(_00030_));
 sky130_fd_sc_hd__o21ai_1 _06656_ (.A1(_00028_),
    .A2(_00029_),
    .B1(_05723_),
    .Y(_00031_));
 sky130_fd_sc_hd__a21bo_1 _06657_ (.A1(_05625_),
    .A2(_05686_),
    .B1_N(_05685_),
    .X(_00032_));
 sky130_fd_sc_hd__and3_1 _06658_ (.A(_00030_),
    .B(_00031_),
    .C(_00032_),
    .X(_00033_));
 sky130_fd_sc_hd__a21oi_1 _06659_ (.A1(_00030_),
    .A2(_00031_),
    .B1(_00032_),
    .Y(_00034_));
 sky130_fd_sc_hd__nor3_1 _06660_ (.A(_05702_),
    .B(_00033_),
    .C(_00034_),
    .Y(_00035_));
 sky130_fd_sc_hd__o21a_1 _06661_ (.A1(_00033_),
    .A2(_00034_),
    .B1(_05702_),
    .X(_00036_));
 sky130_fd_sc_hd__nor2_1 _06662_ (.A(_00035_),
    .B(_00036_),
    .Y(_00037_));
 sky130_fd_sc_hd__and2b_1 _06663_ (.A_N(_05701_),
    .B(_00037_),
    .X(_00038_));
 sky130_fd_sc_hd__xnor2_1 _06664_ (.A(_05701_),
    .B(_00037_),
    .Y(_00039_));
 sky130_fd_sc_hd__and2b_1 _06665_ (.A_N(_05694_),
    .B(_00039_),
    .X(_00040_));
 sky130_fd_sc_hd__xnor2_1 _06666_ (.A(_05694_),
    .B(_00039_),
    .Y(_00041_));
 sky130_fd_sc_hd__and2_1 _06667_ (.A(_05696_),
    .B(_00041_),
    .X(_00042_));
 sky130_fd_sc_hd__nor2_1 _06668_ (.A(_05696_),
    .B(_00041_),
    .Y(_00043_));
 sky130_fd_sc_hd__nor2_1 _06669_ (.A(_00042_),
    .B(_00043_),
    .Y(_00044_));
 sky130_fd_sc_hd__o21ai_1 _06670_ (.A1(_05520_),
    .A2(_05698_),
    .B1(_05604_),
    .Y(_00045_));
 sky130_fd_sc_hd__o21ai_1 _06671_ (.A1(_05525_),
    .A2(_00045_),
    .B1(_05699_),
    .Y(_00046_));
 sky130_fd_sc_hd__and2_1 _06672_ (.A(_05608_),
    .B(_05698_),
    .X(_00047_));
 sky130_fd_sc_hd__a21oi_1 _06673_ (.A1(_05524_),
    .A2(_00047_),
    .B1(_00046_),
    .Y(_00048_));
 sky130_fd_sc_hd__and2b_1 _06674_ (.A_N(_00048_),
    .B(_00044_),
    .X(_00049_));
 sky130_fd_sc_hd__and2b_1 _06675_ (.A_N(_00044_),
    .B(_00048_),
    .X(_00050_));
 sky130_fd_sc_hd__nor2_1 _06676_ (.A(_00049_),
    .B(_00050_),
    .Y(net74));
 sky130_fd_sc_hd__a21o_1 _06677_ (.A1(_05703_),
    .A2(_05722_),
    .B1(_05721_),
    .X(_00051_));
 sky130_fd_sc_hd__o21ba_1 _06678_ (.A1(_05715_),
    .A2(_05716_),
    .B1_N(_05719_),
    .X(_00052_));
 sky130_fd_sc_hd__a22o_1 _06679_ (.A1(net12),
    .A2(net42),
    .B1(net43),
    .B2(net1),
    .X(_00053_));
 sky130_fd_sc_hd__nand2_1 _06680_ (.A(net12),
    .B(net43),
    .Y(_00054_));
 sky130_fd_sc_hd__nor2_1 _06681_ (.A(_05718_),
    .B(_00054_),
    .Y(_00055_));
 sky130_fd_sc_hd__or2_1 _06682_ (.A(_05718_),
    .B(_00054_),
    .X(_00056_));
 sky130_fd_sc_hd__a31o_1 _06683_ (.A1(net12),
    .A2(net41),
    .A3(_05709_),
    .B1(_05707_),
    .X(_00057_));
 sky130_fd_sc_hd__o21ba_1 _06684_ (.A1(_05725_),
    .A2(_05727_),
    .B1_N(_05726_),
    .X(_00058_));
 sky130_fd_sc_hd__and4_1 _06685_ (.A(net27),
    .B(net26),
    .C(net39),
    .D(net40),
    .X(_00059_));
 sky130_fd_sc_hd__a22oi_1 _06686_ (.A1(net27),
    .A2(net39),
    .B1(net40),
    .B2(net26),
    .Y(_00060_));
 sky130_fd_sc_hd__nor2_1 _06687_ (.A(_00059_),
    .B(_00060_),
    .Y(_00061_));
 sky130_fd_sc_hd__nand2_1 _06688_ (.A(net23),
    .B(net41),
    .Y(_00062_));
 sky130_fd_sc_hd__xnor2_1 _06689_ (.A(_00061_),
    .B(_00062_),
    .Y(_00063_));
 sky130_fd_sc_hd__nand2b_1 _06690_ (.A_N(_00058_),
    .B(_00063_),
    .Y(_00064_));
 sky130_fd_sc_hd__xnor2_1 _06691_ (.A(_00058_),
    .B(_00063_),
    .Y(_00065_));
 sky130_fd_sc_hd__nand2_1 _06692_ (.A(_00057_),
    .B(_00065_),
    .Y(_00066_));
 sky130_fd_sc_hd__xnor2_1 _06693_ (.A(_00057_),
    .B(_00065_),
    .Y(_00067_));
 sky130_fd_sc_hd__a21o_1 _06694_ (.A1(_05712_),
    .A2(_05714_),
    .B1(_00067_),
    .X(_00068_));
 sky130_fd_sc_hd__nand3_1 _06695_ (.A(_05712_),
    .B(_05714_),
    .C(_00067_),
    .Y(_00069_));
 sky130_fd_sc_hd__and4_1 _06696_ (.A(_00053_),
    .B(_00056_),
    .C(_00068_),
    .D(_00069_),
    .X(_00070_));
 sky130_fd_sc_hd__nand4_1 _06697_ (.A(_00053_),
    .B(_00056_),
    .C(_00068_),
    .D(_00069_),
    .Y(_00071_));
 sky130_fd_sc_hd__a22oi_1 _06698_ (.A1(_00053_),
    .A2(_00056_),
    .B1(_00068_),
    .B2(_00069_),
    .Y(_00072_));
 sky130_fd_sc_hd__a211oi_1 _06699_ (.A1(_05740_),
    .A2(_05743_),
    .B1(_00070_),
    .C1(_00072_),
    .Y(_00073_));
 sky130_fd_sc_hd__o211a_1 _06700_ (.A1(_00070_),
    .A2(_00072_),
    .B1(_05740_),
    .C1(_05743_),
    .X(_00074_));
 sky130_fd_sc_hd__nor3_1 _06701_ (.A(_00052_),
    .B(_00073_),
    .C(_00074_),
    .Y(_00075_));
 sky130_fd_sc_hd__o21a_1 _06702_ (.A1(_00073_),
    .A2(_00074_),
    .B1(_00052_),
    .X(_00076_));
 sky130_fd_sc_hd__nand2_1 _06703_ (.A(net28),
    .B(net38),
    .Y(_00077_));
 sky130_fd_sc_hd__and4_1 _06704_ (.A(net29),
    .B(net30),
    .C(net36),
    .D(net37),
    .X(_00078_));
 sky130_fd_sc_hd__a22oi_1 _06705_ (.A1(net30),
    .A2(net36),
    .B1(net37),
    .B2(net29),
    .Y(_00079_));
 sky130_fd_sc_hd__nor2_1 _06706_ (.A(_00078_),
    .B(_00079_),
    .Y(_00080_));
 sky130_fd_sc_hd__xnor2_1 _06707_ (.A(_00077_),
    .B(_00080_),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_1 _06708_ (.A(net31),
    .B(net35),
    .Y(_00082_));
 sky130_fd_sc_hd__and4_1 _06709_ (.A(net2),
    .B(net32),
    .C(net64),
    .D(net34),
    .X(_00083_));
 sky130_fd_sc_hd__a22oi_1 _06710_ (.A1(net2),
    .A2(net64),
    .B1(net34),
    .B2(net32),
    .Y(_00084_));
 sky130_fd_sc_hd__nor2_1 _06711_ (.A(_00083_),
    .B(_00084_),
    .Y(_00085_));
 sky130_fd_sc_hd__xnor2_1 _06712_ (.A(_00082_),
    .B(_00085_),
    .Y(_00086_));
 sky130_fd_sc_hd__o21ba_1 _06713_ (.A1(_05730_),
    .A2(_05732_),
    .B1_N(_05731_),
    .X(_00087_));
 sky130_fd_sc_hd__and2b_1 _06714_ (.A_N(_00087_),
    .B(_00086_),
    .X(_00088_));
 sky130_fd_sc_hd__xnor2_1 _06715_ (.A(_00086_),
    .B(_00087_),
    .Y(_00089_));
 sky130_fd_sc_hd__and2_1 _06716_ (.A(_00081_),
    .B(_00089_),
    .X(_00090_));
 sky130_fd_sc_hd__xnor2_1 _06717_ (.A(_00081_),
    .B(_00089_),
    .Y(_00091_));
 sky130_fd_sc_hd__a21o_2 _06718_ (.A1(_05752_),
    .A2(_00000_),
    .B1(_00091_),
    .X(_00092_));
 sky130_fd_sc_hd__nand3_2 _06719_ (.A(_05752_),
    .B(_00000_),
    .C(_00091_),
    .Y(_00093_));
 sky130_fd_sc_hd__o211a_1 _06720_ (.A1(_05736_),
    .A2(_05738_),
    .B1(_00092_),
    .C1(_00093_),
    .X(_00094_));
 sky130_fd_sc_hd__o211ai_2 _06721_ (.A1(_05736_),
    .A2(_05738_),
    .B1(_00092_),
    .C1(_00093_),
    .Y(_00095_));
 sky130_fd_sc_hd__a211oi_2 _06722_ (.A1(_00092_),
    .A2(_00093_),
    .B1(_05736_),
    .C1(_05738_),
    .Y(_00096_));
 sky130_fd_sc_hd__o21ba_1 _06723_ (.A1(_05747_),
    .A2(_05749_),
    .B1_N(_05748_),
    .X(_00097_));
 sky130_fd_sc_hd__o21ba_1 _06724_ (.A1(_00002_),
    .A2(_00004_),
    .B1_N(_00003_),
    .X(_00098_));
 sky130_fd_sc_hd__nand2_1 _06725_ (.A(net63),
    .B(net3),
    .Y(_00099_));
 sky130_fd_sc_hd__and4_1 _06726_ (.A(net61),
    .B(net62),
    .C(net4),
    .D(net5),
    .X(_00100_));
 sky130_fd_sc_hd__a22oi_1 _06727_ (.A1(net62),
    .A2(net4),
    .B1(net5),
    .B2(net61),
    .Y(_00101_));
 sky130_fd_sc_hd__nor2_1 _06728_ (.A(_00100_),
    .B(_00101_),
    .Y(_00102_));
 sky130_fd_sc_hd__xnor2_1 _06729_ (.A(_00099_),
    .B(_00102_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2b_1 _06730_ (.A_N(_00098_),
    .B(_00103_),
    .Y(_00104_));
 sky130_fd_sc_hd__xnor2_1 _06731_ (.A(_00098_),
    .B(_00103_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand2b_1 _06732_ (.A_N(_00097_),
    .B(_00105_),
    .Y(_00106_));
 sky130_fd_sc_hd__xnor2_1 _06733_ (.A(_00097_),
    .B(_00105_),
    .Y(_00107_));
 sky130_fd_sc_hd__nand2_1 _06734_ (.A(net60),
    .B(net6),
    .Y(_00108_));
 sky130_fd_sc_hd__and4_1 _06735_ (.A(net58),
    .B(net59),
    .C(net7),
    .D(net8),
    .X(_00109_));
 sky130_fd_sc_hd__a22oi_1 _06736_ (.A1(net59),
    .A2(net7),
    .B1(net8),
    .B2(net58),
    .Y(_00110_));
 sky130_fd_sc_hd__nor2_1 _06737_ (.A(_00109_),
    .B(_00110_),
    .Y(_00111_));
 sky130_fd_sc_hd__xnor2_1 _06738_ (.A(_00108_),
    .B(_00111_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_1 _06739_ (.A(net55),
    .B(net9),
    .Y(_00113_));
 sky130_fd_sc_hd__and4_1 _06740_ (.A(net33),
    .B(net44),
    .C(net10),
    .D(net11),
    .X(_00114_));
 sky130_fd_sc_hd__a22oi_2 _06741_ (.A1(net44),
    .A2(net10),
    .B1(net11),
    .B2(net33),
    .Y(_00115_));
 sky130_fd_sc_hd__or3_1 _06742_ (.A(_00113_),
    .B(_00114_),
    .C(_00115_),
    .X(_00116_));
 sky130_fd_sc_hd__o21ai_1 _06743_ (.A1(_00114_),
    .A2(_00115_),
    .B1(_00113_),
    .Y(_00117_));
 sky130_fd_sc_hd__o21bai_1 _06744_ (.A1(_00007_),
    .A2(_00009_),
    .B1_N(_00008_),
    .Y(_00118_));
 sky130_fd_sc_hd__nand3_1 _06745_ (.A(_00116_),
    .B(_00117_),
    .C(_00118_),
    .Y(_00119_));
 sky130_fd_sc_hd__a21o_1 _06746_ (.A1(_00116_),
    .A2(_00117_),
    .B1(_00118_),
    .X(_00120_));
 sky130_fd_sc_hd__nand3_1 _06747_ (.A(_00112_),
    .B(_00119_),
    .C(_00120_),
    .Y(_00121_));
 sky130_fd_sc_hd__a21o_1 _06748_ (.A1(_00119_),
    .A2(_00120_),
    .B1(_00112_),
    .X(_00122_));
 sky130_fd_sc_hd__a21bo_1 _06749_ (.A1(_00006_),
    .A2(_00014_),
    .B1_N(_00013_),
    .X(_00123_));
 sky130_fd_sc_hd__nand3_4 _06750_ (.A(_00121_),
    .B(_00122_),
    .C(_00123_),
    .Y(_00124_));
 sky130_fd_sc_hd__a21o_1 _06751_ (.A1(_00121_),
    .A2(_00122_),
    .B1(_00123_),
    .X(_00125_));
 sky130_fd_sc_hd__and3_1 _06752_ (.A(_00107_),
    .B(_00124_),
    .C(_00125_),
    .X(_00126_));
 sky130_fd_sc_hd__nand3_2 _06753_ (.A(_00107_),
    .B(_00124_),
    .C(_00125_),
    .Y(_00127_));
 sky130_fd_sc_hd__a21oi_2 _06754_ (.A1(_00124_),
    .A2(_00125_),
    .B1(_00107_),
    .Y(_00128_));
 sky130_fd_sc_hd__a211oi_4 _06755_ (.A1(_00018_),
    .A2(_00021_),
    .B1(_00126_),
    .C1(_00128_),
    .Y(_00129_));
 sky130_fd_sc_hd__o211a_1 _06756_ (.A1(_00126_),
    .A2(_00128_),
    .B1(_00018_),
    .C1(_00021_),
    .X(_00130_));
 sky130_fd_sc_hd__nor4_2 _06757_ (.A(_00094_),
    .B(_00096_),
    .C(_00129_),
    .D(_00130_),
    .Y(_00131_));
 sky130_fd_sc_hd__or4_1 _06758_ (.A(_00094_),
    .B(_00096_),
    .C(_00129_),
    .D(_00130_),
    .X(_00132_));
 sky130_fd_sc_hd__o22ai_2 _06759_ (.A1(_00094_),
    .A2(_00096_),
    .B1(_00129_),
    .B2(_00130_),
    .Y(_00133_));
 sky130_fd_sc_hd__o211ai_2 _06760_ (.A1(_00023_),
    .A2(_00025_),
    .B1(_00132_),
    .C1(_00133_),
    .Y(_00134_));
 sky130_fd_sc_hd__a211o_1 _06761_ (.A1(_00132_),
    .A2(_00133_),
    .B1(_00023_),
    .C1(_00025_),
    .X(_00135_));
 sky130_fd_sc_hd__or4bb_2 _06762_ (.A(_00075_),
    .B(_00076_),
    .C_N(_00134_),
    .D_N(_00135_),
    .X(_00136_));
 sky130_fd_sc_hd__a2bb2o_1 _06763_ (.A1_N(_00075_),
    .A2_N(_00076_),
    .B1(_00134_),
    .B2(_00135_),
    .X(_00137_));
 sky130_fd_sc_hd__nand2_1 _06764_ (.A(_00136_),
    .B(_00137_),
    .Y(_00138_));
 sky130_fd_sc_hd__nand2b_1 _06765_ (.A_N(_00028_),
    .B(_00030_),
    .Y(_00139_));
 sky130_fd_sc_hd__xnor2_1 _06766_ (.A(_00138_),
    .B(_00139_),
    .Y(_00140_));
 sky130_fd_sc_hd__xnor2_1 _06767_ (.A(_00051_),
    .B(_00140_),
    .Y(_00141_));
 sky130_fd_sc_hd__nor2_1 _06768_ (.A(_00033_),
    .B(_00035_),
    .Y(_00142_));
 sky130_fd_sc_hd__or2_1 _06769_ (.A(_00141_),
    .B(_00142_),
    .X(_00143_));
 sky130_fd_sc_hd__xor2_1 _06770_ (.A(_00141_),
    .B(_00142_),
    .X(_00144_));
 sky130_fd_sc_hd__and2_1 _06771_ (.A(_00038_),
    .B(_00144_),
    .X(_00145_));
 sky130_fd_sc_hd__nor2_1 _06772_ (.A(_00038_),
    .B(_00144_),
    .Y(_00146_));
 sky130_fd_sc_hd__nor2_1 _06773_ (.A(_00145_),
    .B(_00146_),
    .Y(_00147_));
 sky130_fd_sc_hd__xor2_1 _06774_ (.A(_00040_),
    .B(_00147_),
    .X(_00148_));
 sky130_fd_sc_hd__nor2_1 _06775_ (.A(_00042_),
    .B(_00049_),
    .Y(_00149_));
 sky130_fd_sc_hd__xnor2_1 _06776_ (.A(_00148_),
    .B(_00149_),
    .Y(net75));
 sky130_fd_sc_hd__nor2_1 _06777_ (.A(_00073_),
    .B(_00075_),
    .Y(_00150_));
 sky130_fd_sc_hd__and4_1 _06778_ (.A(net23),
    .B(net12),
    .C(net42),
    .D(net43),
    .X(_00151_));
 sky130_fd_sc_hd__nand2_1 _06779_ (.A(net23),
    .B(net42),
    .Y(_00152_));
 sky130_fd_sc_hd__a21oi_1 _06780_ (.A1(_00054_),
    .A2(_00152_),
    .B1(_00151_),
    .Y(_00153_));
 sky130_fd_sc_hd__nand2_1 _06781_ (.A(net1),
    .B(net45),
    .Y(_00154_));
 sky130_fd_sc_hd__xnor2_1 _06782_ (.A(_00153_),
    .B(_00154_),
    .Y(_00155_));
 sky130_fd_sc_hd__and2_1 _06783_ (.A(_00055_),
    .B(_00155_),
    .X(_00156_));
 sky130_fd_sc_hd__nor2_1 _06784_ (.A(_00055_),
    .B(_00155_),
    .Y(_00157_));
 sky130_fd_sc_hd__or2_1 _06785_ (.A(_00156_),
    .B(_00157_),
    .X(_00158_));
 sky130_fd_sc_hd__a31o_1 _06786_ (.A1(net23),
    .A2(net41),
    .A3(_00061_),
    .B1(_00059_),
    .X(_00159_));
 sky130_fd_sc_hd__o21ba_1 _06787_ (.A1(_00077_),
    .A2(_00079_),
    .B1_N(_00078_),
    .X(_00160_));
 sky130_fd_sc_hd__and4_1 _06788_ (.A(net28),
    .B(net27),
    .C(net39),
    .D(net40),
    .X(_00161_));
 sky130_fd_sc_hd__a22oi_1 _06789_ (.A1(net28),
    .A2(net39),
    .B1(net40),
    .B2(net27),
    .Y(_00162_));
 sky130_fd_sc_hd__nor2_1 _06790_ (.A(_00161_),
    .B(_00162_),
    .Y(_00163_));
 sky130_fd_sc_hd__nand2_1 _06791_ (.A(net26),
    .B(net41),
    .Y(_00164_));
 sky130_fd_sc_hd__xnor2_1 _06792_ (.A(_00163_),
    .B(_00164_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2b_1 _06793_ (.A_N(_00160_),
    .B(_00165_),
    .Y(_00166_));
 sky130_fd_sc_hd__xnor2_1 _06794_ (.A(_00160_),
    .B(_00165_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand2_1 _06795_ (.A(_00159_),
    .B(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__xnor2_1 _06796_ (.A(_00159_),
    .B(_00167_),
    .Y(_00169_));
 sky130_fd_sc_hd__a21oi_2 _06797_ (.A1(_00064_),
    .A2(_00066_),
    .B1(_00169_),
    .Y(_00170_));
 sky130_fd_sc_hd__inv_2 _06798_ (.A(_00170_),
    .Y(_00171_));
 sky130_fd_sc_hd__and3_1 _06799_ (.A(_00064_),
    .B(_00066_),
    .C(_00169_),
    .X(_00172_));
 sky130_fd_sc_hd__nor3_1 _06800_ (.A(_00158_),
    .B(_00170_),
    .C(_00172_),
    .Y(_00173_));
 sky130_fd_sc_hd__or3_1 _06801_ (.A(_00158_),
    .B(_00170_),
    .C(_00172_),
    .X(_00174_));
 sky130_fd_sc_hd__o21a_1 _06802_ (.A1(_00170_),
    .A2(_00172_),
    .B1(_00158_),
    .X(_00175_));
 sky130_fd_sc_hd__a211oi_2 _06803_ (.A1(_00092_),
    .A2(_00095_),
    .B1(_00173_),
    .C1(_00175_),
    .Y(_00176_));
 sky130_fd_sc_hd__o211a_1 _06804_ (.A1(_00173_),
    .A2(_00175_),
    .B1(_00092_),
    .C1(_00095_),
    .X(_00177_));
 sky130_fd_sc_hd__a211oi_2 _06805_ (.A1(_00068_),
    .A2(_00071_),
    .B1(_00176_),
    .C1(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__o211a_1 _06806_ (.A1(_00176_),
    .A2(_00177_),
    .B1(_00068_),
    .C1(_00071_),
    .X(_00179_));
 sky130_fd_sc_hd__nand2_1 _06807_ (.A(net29),
    .B(net38),
    .Y(_00180_));
 sky130_fd_sc_hd__and4_1 _06808_ (.A(net30),
    .B(net31),
    .C(net36),
    .D(net37),
    .X(_00181_));
 sky130_fd_sc_hd__a22oi_1 _06809_ (.A1(net31),
    .A2(net36),
    .B1(net37),
    .B2(net30),
    .Y(_00182_));
 sky130_fd_sc_hd__nor2_1 _06810_ (.A(_00181_),
    .B(_00182_),
    .Y(_00183_));
 sky130_fd_sc_hd__xnor2_1 _06811_ (.A(_00180_),
    .B(_00183_),
    .Y(_00184_));
 sky130_fd_sc_hd__nand2_1 _06812_ (.A(net32),
    .B(net35),
    .Y(_00185_));
 sky130_fd_sc_hd__and4_1 _06813_ (.A(net2),
    .B(net64),
    .C(net34),
    .D(net3),
    .X(_00186_));
 sky130_fd_sc_hd__a22oi_1 _06814_ (.A1(net2),
    .A2(net34),
    .B1(net3),
    .B2(net64),
    .Y(_00187_));
 sky130_fd_sc_hd__nor2_1 _06815_ (.A(_00186_),
    .B(_00187_),
    .Y(_00188_));
 sky130_fd_sc_hd__xnor2_1 _06816_ (.A(_00185_),
    .B(_00188_),
    .Y(_00189_));
 sky130_fd_sc_hd__o21ba_1 _06817_ (.A1(_00082_),
    .A2(_00084_),
    .B1_N(_00083_),
    .X(_00190_));
 sky130_fd_sc_hd__and2b_1 _06818_ (.A_N(_00190_),
    .B(_00189_),
    .X(_00191_));
 sky130_fd_sc_hd__xnor2_1 _06819_ (.A(_00189_),
    .B(_00190_),
    .Y(_00192_));
 sky130_fd_sc_hd__and2_1 _06820_ (.A(_00184_),
    .B(_00192_),
    .X(_00193_));
 sky130_fd_sc_hd__xnor2_1 _06821_ (.A(_00184_),
    .B(_00192_),
    .Y(_00194_));
 sky130_fd_sc_hd__a21o_2 _06822_ (.A1(_00104_),
    .A2(_00106_),
    .B1(_00194_),
    .X(_00195_));
 sky130_fd_sc_hd__nand3_2 _06823_ (.A(_00104_),
    .B(_00106_),
    .C(_00194_),
    .Y(_00196_));
 sky130_fd_sc_hd__o211a_1 _06824_ (.A1(_00088_),
    .A2(_00090_),
    .B1(_00195_),
    .C1(_00196_),
    .X(_00197_));
 sky130_fd_sc_hd__o211ai_2 _06825_ (.A1(_00088_),
    .A2(_00090_),
    .B1(_00195_),
    .C1(_00196_),
    .Y(_00198_));
 sky130_fd_sc_hd__a211oi_2 _06826_ (.A1(_00195_),
    .A2(_00196_),
    .B1(_00088_),
    .C1(_00090_),
    .Y(_00199_));
 sky130_fd_sc_hd__o21ba_1 _06827_ (.A1(_00099_),
    .A2(_00101_),
    .B1_N(_00100_),
    .X(_00200_));
 sky130_fd_sc_hd__o21ba_1 _06828_ (.A1(_00108_),
    .A2(_00110_),
    .B1_N(_00109_),
    .X(_00201_));
 sky130_fd_sc_hd__and4_1 _06829_ (.A(net61),
    .B(net62),
    .C(net5),
    .D(net6),
    .X(_00202_));
 sky130_fd_sc_hd__a22oi_1 _06830_ (.A1(net62),
    .A2(net5),
    .B1(net6),
    .B2(net61),
    .Y(_00203_));
 sky130_fd_sc_hd__nor2_1 _06831_ (.A(_00202_),
    .B(_00203_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _06832_ (.A(net63),
    .B(net4),
    .Y(_00205_));
 sky130_fd_sc_hd__xnor2_1 _06833_ (.A(_00204_),
    .B(_00205_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2b_1 _06834_ (.A_N(_00201_),
    .B(_00206_),
    .Y(_00207_));
 sky130_fd_sc_hd__xnor2_1 _06835_ (.A(_00201_),
    .B(_00206_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2b_1 _06836_ (.A_N(_00200_),
    .B(_00208_),
    .Y(_00209_));
 sky130_fd_sc_hd__xnor2_1 _06837_ (.A(_00200_),
    .B(_00208_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _06838_ (.A(net60),
    .B(net7),
    .Y(_00211_));
 sky130_fd_sc_hd__and4_1 _06839_ (.A(net58),
    .B(net59),
    .C(net8),
    .D(net9),
    .X(_00212_));
 sky130_fd_sc_hd__a22oi_1 _06840_ (.A1(net59),
    .A2(net8),
    .B1(net9),
    .B2(net58),
    .Y(_00213_));
 sky130_fd_sc_hd__nor2_1 _06841_ (.A(_00212_),
    .B(_00213_),
    .Y(_00214_));
 sky130_fd_sc_hd__xnor2_1 _06842_ (.A(_00211_),
    .B(_00214_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _06843_ (.A(net55),
    .B(net10),
    .Y(_00216_));
 sky130_fd_sc_hd__and4_1 _06844_ (.A(net33),
    .B(net44),
    .C(net11),
    .D(net13),
    .X(_00217_));
 sky130_fd_sc_hd__a22oi_2 _06845_ (.A1(net44),
    .A2(net11),
    .B1(net13),
    .B2(net33),
    .Y(_00218_));
 sky130_fd_sc_hd__or3_1 _06846_ (.A(_00216_),
    .B(_00217_),
    .C(_00218_),
    .X(_00219_));
 sky130_fd_sc_hd__o21ai_1 _06847_ (.A1(_00217_),
    .A2(_00218_),
    .B1(_00216_),
    .Y(_00220_));
 sky130_fd_sc_hd__o21bai_1 _06848_ (.A1(_00113_),
    .A2(_00115_),
    .B1_N(_00114_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand3_1 _06849_ (.A(_00219_),
    .B(_00220_),
    .C(_00221_),
    .Y(_00222_));
 sky130_fd_sc_hd__a21o_1 _06850_ (.A1(_00219_),
    .A2(_00220_),
    .B1(_00221_),
    .X(_00223_));
 sky130_fd_sc_hd__nand3_1 _06851_ (.A(_00215_),
    .B(_00222_),
    .C(_00223_),
    .Y(_00224_));
 sky130_fd_sc_hd__a21o_1 _06852_ (.A1(_00222_),
    .A2(_00223_),
    .B1(_00215_),
    .X(_00225_));
 sky130_fd_sc_hd__a21bo_1 _06853_ (.A1(_00112_),
    .A2(_00120_),
    .B1_N(_00119_),
    .X(_00226_));
 sky130_fd_sc_hd__nand3_4 _06854_ (.A(_00224_),
    .B(_00225_),
    .C(_00226_),
    .Y(_00227_));
 sky130_fd_sc_hd__a21o_1 _06855_ (.A1(_00224_),
    .A2(_00225_),
    .B1(_00226_),
    .X(_00228_));
 sky130_fd_sc_hd__and3_1 _06856_ (.A(_00210_),
    .B(_00227_),
    .C(_00228_),
    .X(_00229_));
 sky130_fd_sc_hd__nand3_2 _06857_ (.A(_00210_),
    .B(_00227_),
    .C(_00228_),
    .Y(_00230_));
 sky130_fd_sc_hd__a21oi_2 _06858_ (.A1(_00227_),
    .A2(_00228_),
    .B1(_00210_),
    .Y(_00231_));
 sky130_fd_sc_hd__a211oi_4 _06859_ (.A1(_00124_),
    .A2(_00127_),
    .B1(_00229_),
    .C1(_00231_),
    .Y(_00232_));
 sky130_fd_sc_hd__o211a_1 _06860_ (.A1(_00229_),
    .A2(_00231_),
    .B1(_00124_),
    .C1(_00127_),
    .X(_00233_));
 sky130_fd_sc_hd__nor4_2 _06861_ (.A(_00197_),
    .B(_00199_),
    .C(_00232_),
    .D(_00233_),
    .Y(_00234_));
 sky130_fd_sc_hd__or4_2 _06862_ (.A(_00197_),
    .B(_00199_),
    .C(_00232_),
    .D(_00233_),
    .X(_00235_));
 sky130_fd_sc_hd__o22ai_2 _06863_ (.A1(_00197_),
    .A2(_00199_),
    .B1(_00232_),
    .B2(_00233_),
    .Y(_00236_));
 sky130_fd_sc_hd__o211ai_4 _06864_ (.A1(_00129_),
    .A2(_00131_),
    .B1(_00235_),
    .C1(_00236_),
    .Y(_00237_));
 sky130_fd_sc_hd__a211o_1 _06865_ (.A1(_00235_),
    .A2(_00236_),
    .B1(_00129_),
    .C1(_00131_),
    .X(_00238_));
 sky130_fd_sc_hd__and4bb_1 _06866_ (.A_N(_00178_),
    .B_N(_00179_),
    .C(_00237_),
    .D(_00238_),
    .X(_00239_));
 sky130_fd_sc_hd__or4bb_1 _06867_ (.A(_00178_),
    .B(_00179_),
    .C_N(_00237_),
    .D_N(_00238_),
    .X(_00240_));
 sky130_fd_sc_hd__a2bb2oi_1 _06868_ (.A1_N(_00178_),
    .A2_N(_00179_),
    .B1(_00237_),
    .B2(_00238_),
    .Y(_00241_));
 sky130_fd_sc_hd__a211oi_2 _06869_ (.A1(_00134_),
    .A2(_00136_),
    .B1(_00239_),
    .C1(_00241_),
    .Y(_00242_));
 sky130_fd_sc_hd__o211a_1 _06870_ (.A1(_00239_),
    .A2(_00241_),
    .B1(_00134_),
    .C1(_00136_),
    .X(_00243_));
 sky130_fd_sc_hd__nor2_1 _06871_ (.A(_00242_),
    .B(_00243_),
    .Y(_00244_));
 sky130_fd_sc_hd__and2b_1 _06872_ (.A_N(_00150_),
    .B(_00244_),
    .X(_00245_));
 sky130_fd_sc_hd__xnor2_1 _06873_ (.A(_00150_),
    .B(_00244_),
    .Y(_00246_));
 sky130_fd_sc_hd__a32oi_2 _06874_ (.A1(_00136_),
    .A2(_00137_),
    .A3(_00139_),
    .B1(_00140_),
    .B2(_00051_),
    .Y(_00247_));
 sky130_fd_sc_hd__and2b_1 _06875_ (.A_N(_00247_),
    .B(_00246_),
    .X(_00248_));
 sky130_fd_sc_hd__xnor2_1 _06876_ (.A(_00246_),
    .B(_00247_),
    .Y(_00249_));
 sky130_fd_sc_hd__and2b_1 _06877_ (.A_N(_00143_),
    .B(_00249_),
    .X(_00250_));
 sky130_fd_sc_hd__xnor2_1 _06878_ (.A(_00143_),
    .B(_00249_),
    .Y(_00251_));
 sky130_fd_sc_hd__and2_1 _06879_ (.A(_00145_),
    .B(_00251_),
    .X(_00252_));
 sky130_fd_sc_hd__xor2_1 _06880_ (.A(_00145_),
    .B(_00251_),
    .X(_00253_));
 sky130_fd_sc_hd__inv_2 _06881_ (.A(_00253_),
    .Y(_00254_));
 sky130_fd_sc_hd__and2_1 _06882_ (.A(_00044_),
    .B(_00148_),
    .X(_00255_));
 sky130_fd_sc_hd__o21a_1 _06883_ (.A1(_00040_),
    .A2(_00042_),
    .B1(_00147_),
    .X(_00256_));
 sky130_fd_sc_hd__a31o_1 _06884_ (.A1(_00044_),
    .A2(_00046_),
    .A3(_00148_),
    .B1(_00256_),
    .X(_00257_));
 sky130_fd_sc_hd__a31oi_2 _06885_ (.A1(_05524_),
    .A2(_00047_),
    .A3(_00255_),
    .B1(_00257_),
    .Y(_00258_));
 sky130_fd_sc_hd__nor2_1 _06886_ (.A(_00254_),
    .B(_00258_),
    .Y(_00259_));
 sky130_fd_sc_hd__xnor2_1 _06887_ (.A(_00253_),
    .B(_00258_),
    .Y(net77));
 sky130_fd_sc_hd__o21ai_1 _06888_ (.A1(_00176_),
    .A2(_00178_),
    .B1(_00156_),
    .Y(_00260_));
 sky130_fd_sc_hd__or3_1 _06889_ (.A(_00156_),
    .B(_00176_),
    .C(_00178_),
    .X(_00261_));
 sky130_fd_sc_hd__and2_1 _06890_ (.A(_00260_),
    .B(_00261_),
    .X(_00262_));
 sky130_fd_sc_hd__and4_1 _06891_ (.A(net26),
    .B(net23),
    .C(net42),
    .D(net43),
    .X(_00263_));
 sky130_fd_sc_hd__a22o_1 _06892_ (.A1(net26),
    .A2(net42),
    .B1(net43),
    .B2(net23),
    .X(_00264_));
 sky130_fd_sc_hd__and2b_1 _06893_ (.A_N(_00263_),
    .B(_00264_),
    .X(_00265_));
 sky130_fd_sc_hd__nand2_1 _06894_ (.A(net12),
    .B(net45),
    .Y(_00266_));
 sky130_fd_sc_hd__xnor2_1 _06895_ (.A(_00265_),
    .B(_00266_),
    .Y(_00267_));
 sky130_fd_sc_hd__a31oi_1 _06896_ (.A1(net1),
    .A2(net45),
    .A3(_00153_),
    .B1(_00151_),
    .Y(_00268_));
 sky130_fd_sc_hd__and2b_1 _06897_ (.A_N(_00268_),
    .B(_00267_),
    .X(_00269_));
 sky130_fd_sc_hd__xnor2_1 _06898_ (.A(_00267_),
    .B(_00268_),
    .Y(_00270_));
 sky130_fd_sc_hd__nand2_1 _06899_ (.A(net1),
    .B(net46),
    .Y(_00271_));
 sky130_fd_sc_hd__xor2_1 _06900_ (.A(_00270_),
    .B(_00271_),
    .X(_00272_));
 sky130_fd_sc_hd__a31o_1 _06901_ (.A1(net26),
    .A2(net41),
    .A3(_00163_),
    .B1(_00161_),
    .X(_00273_));
 sky130_fd_sc_hd__o21ba_1 _06902_ (.A1(_00180_),
    .A2(_00182_),
    .B1_N(_00181_),
    .X(_00274_));
 sky130_fd_sc_hd__and4_1 _06903_ (.A(net28),
    .B(net29),
    .C(net39),
    .D(net40),
    .X(_00275_));
 sky130_fd_sc_hd__a22oi_1 _06904_ (.A1(net29),
    .A2(net39),
    .B1(net40),
    .B2(net28),
    .Y(_00276_));
 sky130_fd_sc_hd__nor2_1 _06905_ (.A(_00275_),
    .B(_00276_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _06906_ (.A(net27),
    .B(net41),
    .Y(_00278_));
 sky130_fd_sc_hd__xnor2_1 _06907_ (.A(_00277_),
    .B(_00278_),
    .Y(_00279_));
 sky130_fd_sc_hd__nand2b_1 _06908_ (.A_N(_00274_),
    .B(_00279_),
    .Y(_00280_));
 sky130_fd_sc_hd__xnor2_1 _06909_ (.A(_00274_),
    .B(_00279_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_1 _06910_ (.A(_00273_),
    .B(_00281_),
    .Y(_00282_));
 sky130_fd_sc_hd__xnor2_1 _06911_ (.A(_00273_),
    .B(_00281_),
    .Y(_00283_));
 sky130_fd_sc_hd__a21oi_2 _06912_ (.A1(_00166_),
    .A2(_00168_),
    .B1(_00283_),
    .Y(_00284_));
 sky130_fd_sc_hd__inv_2 _06913_ (.A(_00284_),
    .Y(_00285_));
 sky130_fd_sc_hd__and3_1 _06914_ (.A(_00166_),
    .B(_00168_),
    .C(_00283_),
    .X(_00286_));
 sky130_fd_sc_hd__nor3_1 _06915_ (.A(_00272_),
    .B(_00284_),
    .C(_00286_),
    .Y(_00288_));
 sky130_fd_sc_hd__or3_1 _06916_ (.A(_00272_),
    .B(_00284_),
    .C(_00286_),
    .X(_00289_));
 sky130_fd_sc_hd__o21a_1 _06917_ (.A1(_00284_),
    .A2(_00286_),
    .B1(_00272_),
    .X(_00290_));
 sky130_fd_sc_hd__a211oi_2 _06918_ (.A1(_00195_),
    .A2(_00198_),
    .B1(_00288_),
    .C1(_00290_),
    .Y(_00291_));
 sky130_fd_sc_hd__o211a_1 _06919_ (.A1(_00288_),
    .A2(_00290_),
    .B1(_00195_),
    .C1(_00198_),
    .X(_00292_));
 sky130_fd_sc_hd__a211oi_2 _06920_ (.A1(_00171_),
    .A2(_00174_),
    .B1(_00291_),
    .C1(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__o211a_1 _06921_ (.A1(_00291_),
    .A2(_00292_),
    .B1(_00171_),
    .C1(_00174_),
    .X(_00294_));
 sky130_fd_sc_hd__and4_1 _06922_ (.A(net31),
    .B(net32),
    .C(net36),
    .D(net37),
    .X(_00295_));
 sky130_fd_sc_hd__a22oi_1 _06923_ (.A1(net32),
    .A2(net36),
    .B1(net37),
    .B2(net31),
    .Y(_00296_));
 sky130_fd_sc_hd__nor2_1 _06924_ (.A(_00295_),
    .B(_00296_),
    .Y(_00297_));
 sky130_fd_sc_hd__nand2_1 _06925_ (.A(net30),
    .B(net38),
    .Y(_00299_));
 sky130_fd_sc_hd__xnor2_1 _06926_ (.A(_00297_),
    .B(_00299_),
    .Y(_00300_));
 sky130_fd_sc_hd__and4_1 _06927_ (.A(net64),
    .B(net34),
    .C(net3),
    .D(net4),
    .X(_00301_));
 sky130_fd_sc_hd__a22oi_1 _06928_ (.A1(net34),
    .A2(net3),
    .B1(net4),
    .B2(net64),
    .Y(_00302_));
 sky130_fd_sc_hd__nor2_1 _06929_ (.A(_00301_),
    .B(_00302_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _06930_ (.A(net2),
    .B(net35),
    .Y(_00304_));
 sky130_fd_sc_hd__xnor2_1 _06931_ (.A(_00303_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__o21ba_1 _06932_ (.A1(_00185_),
    .A2(_00187_),
    .B1_N(_00186_),
    .X(_00306_));
 sky130_fd_sc_hd__and2b_1 _06933_ (.A_N(_00306_),
    .B(_00305_),
    .X(_00307_));
 sky130_fd_sc_hd__xnor2_1 _06934_ (.A(_00305_),
    .B(_00306_),
    .Y(_00308_));
 sky130_fd_sc_hd__and2_1 _06935_ (.A(_00300_),
    .B(_00308_),
    .X(_00310_));
 sky130_fd_sc_hd__xnor2_1 _06936_ (.A(_00300_),
    .B(_00308_),
    .Y(_00311_));
 sky130_fd_sc_hd__a21o_1 _06937_ (.A1(_00207_),
    .A2(_00209_),
    .B1(_00311_),
    .X(_00312_));
 sky130_fd_sc_hd__inv_2 _06938_ (.A(_00312_),
    .Y(_00313_));
 sky130_fd_sc_hd__nand3_1 _06939_ (.A(_00207_),
    .B(_00209_),
    .C(_00311_),
    .Y(_00314_));
 sky130_fd_sc_hd__o211a_1 _06940_ (.A1(_00191_),
    .A2(_00193_),
    .B1(_00312_),
    .C1(_00314_),
    .X(_00315_));
 sky130_fd_sc_hd__a211oi_2 _06941_ (.A1(_00312_),
    .A2(_00314_),
    .B1(_00191_),
    .C1(_00193_),
    .Y(_00316_));
 sky130_fd_sc_hd__o21ba_1 _06942_ (.A1(_00203_),
    .A2(_00205_),
    .B1_N(_00202_),
    .X(_00317_));
 sky130_fd_sc_hd__o21ba_1 _06943_ (.A1(_00211_),
    .A2(_00213_),
    .B1_N(_00212_),
    .X(_00318_));
 sky130_fd_sc_hd__and4_1 _06944_ (.A(net61),
    .B(net62),
    .C(net6),
    .D(net7),
    .X(_00319_));
 sky130_fd_sc_hd__a22oi_1 _06945_ (.A1(net62),
    .A2(net6),
    .B1(net7),
    .B2(net61),
    .Y(_00321_));
 sky130_fd_sc_hd__nor2_1 _06946_ (.A(_00319_),
    .B(_00321_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(net63),
    .B(net5),
    .Y(_00323_));
 sky130_fd_sc_hd__xnor2_1 _06948_ (.A(_00322_),
    .B(_00323_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2b_1 _06949_ (.A_N(_00318_),
    .B(_00324_),
    .Y(_00325_));
 sky130_fd_sc_hd__xnor2_1 _06950_ (.A(_00318_),
    .B(_00324_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2b_1 _06951_ (.A_N(_00317_),
    .B(_00326_),
    .Y(_00327_));
 sky130_fd_sc_hd__xnor2_1 _06952_ (.A(_00317_),
    .B(_00326_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _06953_ (.A(net60),
    .B(net8),
    .Y(_00329_));
 sky130_fd_sc_hd__and4_1 _06954_ (.A(net58),
    .B(net59),
    .C(net9),
    .D(net10),
    .X(_00330_));
 sky130_fd_sc_hd__a22oi_1 _06955_ (.A1(net59),
    .A2(net9),
    .B1(net10),
    .B2(net58),
    .Y(_00332_));
 sky130_fd_sc_hd__nor2_1 _06956_ (.A(_00330_),
    .B(_00332_),
    .Y(_00333_));
 sky130_fd_sc_hd__xnor2_1 _06957_ (.A(_00329_),
    .B(_00333_),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _06958_ (.A(net55),
    .B(net11),
    .Y(_00335_));
 sky130_fd_sc_hd__and4_1 _06959_ (.A(net33),
    .B(net44),
    .C(net13),
    .D(net14),
    .X(_00336_));
 sky130_fd_sc_hd__a22oi_2 _06960_ (.A1(net44),
    .A2(net13),
    .B1(net14),
    .B2(net33),
    .Y(_00337_));
 sky130_fd_sc_hd__or3_1 _06961_ (.A(_00335_),
    .B(_00336_),
    .C(_00337_),
    .X(_00338_));
 sky130_fd_sc_hd__o21ai_1 _06962_ (.A1(_00336_),
    .A2(_00337_),
    .B1(_00335_),
    .Y(_00339_));
 sky130_fd_sc_hd__o21bai_1 _06963_ (.A1(_00216_),
    .A2(_00218_),
    .B1_N(_00217_),
    .Y(_00340_));
 sky130_fd_sc_hd__nand3_1 _06964_ (.A(_00338_),
    .B(_00339_),
    .C(_00340_),
    .Y(_00341_));
 sky130_fd_sc_hd__a21o_1 _06965_ (.A1(_00338_),
    .A2(_00339_),
    .B1(_00340_),
    .X(_00343_));
 sky130_fd_sc_hd__nand3_2 _06966_ (.A(_00334_),
    .B(_00341_),
    .C(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__a21o_1 _06967_ (.A1(_00341_),
    .A2(_00343_),
    .B1(_00334_),
    .X(_00345_));
 sky130_fd_sc_hd__a21bo_1 _06968_ (.A1(_00215_),
    .A2(_00223_),
    .B1_N(_00222_),
    .X(_00346_));
 sky130_fd_sc_hd__nand3_4 _06969_ (.A(_00344_),
    .B(_00345_),
    .C(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__a21o_1 _06970_ (.A1(_00344_),
    .A2(_00345_),
    .B1(_00346_),
    .X(_00348_));
 sky130_fd_sc_hd__and3_1 _06971_ (.A(_00328_),
    .B(_00347_),
    .C(_00348_),
    .X(_00349_));
 sky130_fd_sc_hd__nand3_2 _06972_ (.A(_00328_),
    .B(_00347_),
    .C(_00348_),
    .Y(_00350_));
 sky130_fd_sc_hd__a21oi_2 _06973_ (.A1(_00347_),
    .A2(_00348_),
    .B1(_00328_),
    .Y(_00351_));
 sky130_fd_sc_hd__a211oi_4 _06974_ (.A1(_00227_),
    .A2(_00230_),
    .B1(_00349_),
    .C1(_00351_),
    .Y(_00352_));
 sky130_fd_sc_hd__o211a_1 _06975_ (.A1(_00349_),
    .A2(_00351_),
    .B1(_00227_),
    .C1(_00230_),
    .X(_00354_));
 sky130_fd_sc_hd__nor4_2 _06976_ (.A(_00315_),
    .B(_00316_),
    .C(_00352_),
    .D(_00354_),
    .Y(_00355_));
 sky130_fd_sc_hd__or4_2 _06977_ (.A(_00315_),
    .B(_00316_),
    .C(_00352_),
    .D(_00354_),
    .X(_00356_));
 sky130_fd_sc_hd__o22ai_2 _06978_ (.A1(_00315_),
    .A2(_00316_),
    .B1(_00352_),
    .B2(_00354_),
    .Y(_00357_));
 sky130_fd_sc_hd__o211ai_4 _06979_ (.A1(_00232_),
    .A2(_00234_),
    .B1(_00356_),
    .C1(_00357_),
    .Y(_00358_));
 sky130_fd_sc_hd__a211o_1 _06980_ (.A1(_00356_),
    .A2(_00357_),
    .B1(_00232_),
    .C1(_00234_),
    .X(_00359_));
 sky130_fd_sc_hd__and4bb_1 _06981_ (.A_N(_00293_),
    .B_N(_00294_),
    .C(_00358_),
    .D(_00359_),
    .X(_00360_));
 sky130_fd_sc_hd__or4bb_1 _06982_ (.A(_00293_),
    .B(_00294_),
    .C_N(_00358_),
    .D_N(_00359_),
    .X(_00361_));
 sky130_fd_sc_hd__a2bb2oi_1 _06983_ (.A1_N(_00293_),
    .A2_N(_00294_),
    .B1(_00358_),
    .B2(_00359_),
    .Y(_00362_));
 sky130_fd_sc_hd__a211o_1 _06984_ (.A1(_00237_),
    .A2(_00240_),
    .B1(_00360_),
    .C1(_00362_),
    .X(_00363_));
 sky130_fd_sc_hd__o211ai_2 _06985_ (.A1(_00360_),
    .A2(_00362_),
    .B1(_00237_),
    .C1(_00240_),
    .Y(_00365_));
 sky130_fd_sc_hd__nand3_2 _06986_ (.A(_00262_),
    .B(_00363_),
    .C(_00365_),
    .Y(_00366_));
 sky130_fd_sc_hd__a21o_1 _06987_ (.A1(_00363_),
    .A2(_00365_),
    .B1(_00262_),
    .X(_00367_));
 sky130_fd_sc_hd__o211ai_2 _06988_ (.A1(_00242_),
    .A2(_00245_),
    .B1(_00366_),
    .C1(_00367_),
    .Y(_00368_));
 sky130_fd_sc_hd__a211o_1 _06989_ (.A1(_00366_),
    .A2(_00367_),
    .B1(_00242_),
    .C1(_00245_),
    .X(_00369_));
 sky130_fd_sc_hd__nand2_1 _06990_ (.A(_00368_),
    .B(_00369_),
    .Y(_00370_));
 sky130_fd_sc_hd__and3_1 _06991_ (.A(_00248_),
    .B(_00368_),
    .C(_00369_),
    .X(_00371_));
 sky130_fd_sc_hd__xnor2_1 _06992_ (.A(_00248_),
    .B(_00370_),
    .Y(_00372_));
 sky130_fd_sc_hd__xor2_1 _06993_ (.A(_00250_),
    .B(_00372_),
    .X(_00373_));
 sky130_fd_sc_hd__nor2_1 _06994_ (.A(_00252_),
    .B(_00259_),
    .Y(_00374_));
 sky130_fd_sc_hd__xnor2_1 _06995_ (.A(_00373_),
    .B(_00374_),
    .Y(net78));
 sky130_fd_sc_hd__a31oi_1 _06996_ (.A1(net1),
    .A2(net46),
    .A3(_00270_),
    .B1(_00269_),
    .Y(_00376_));
 sky130_fd_sc_hd__o21ba_1 _06997_ (.A1(_00291_),
    .A2(_00293_),
    .B1_N(_00376_),
    .X(_00377_));
 sky130_fd_sc_hd__or3b_1 _06998_ (.A(_00291_),
    .B(_00293_),
    .C_N(_00376_),
    .X(_00378_));
 sky130_fd_sc_hd__and2b_1 _06999_ (.A_N(_00377_),
    .B(_00378_),
    .X(_00379_));
 sky130_fd_sc_hd__a22o_1 _07000_ (.A1(net12),
    .A2(net46),
    .B1(net47),
    .B2(net1),
    .X(_00380_));
 sky130_fd_sc_hd__nand4_2 _07001_ (.A(net12),
    .B(net1),
    .C(net46),
    .D(net47),
    .Y(_00381_));
 sky130_fd_sc_hd__and4_1 _07002_ (.A(net27),
    .B(net26),
    .C(net42),
    .D(net43),
    .X(_00382_));
 sky130_fd_sc_hd__a22o_1 _07003_ (.A1(net27),
    .A2(net42),
    .B1(net43),
    .B2(net26),
    .X(_00383_));
 sky130_fd_sc_hd__and2b_1 _07004_ (.A_N(_00382_),
    .B(_00383_),
    .X(_00384_));
 sky130_fd_sc_hd__nand2_1 _07005_ (.A(net23),
    .B(net45),
    .Y(_00386_));
 sky130_fd_sc_hd__xnor2_1 _07006_ (.A(_00384_),
    .B(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__a31o_1 _07007_ (.A1(net12),
    .A2(net45),
    .A3(_00264_),
    .B1(_00263_),
    .X(_00388_));
 sky130_fd_sc_hd__nand2_1 _07008_ (.A(_00387_),
    .B(_00388_),
    .Y(_00389_));
 sky130_fd_sc_hd__or2_1 _07009_ (.A(_00387_),
    .B(_00388_),
    .X(_00390_));
 sky130_fd_sc_hd__nand4_2 _07010_ (.A(_00380_),
    .B(_00381_),
    .C(_00389_),
    .D(_00390_),
    .Y(_00391_));
 sky130_fd_sc_hd__a22o_1 _07011_ (.A1(_00380_),
    .A2(_00381_),
    .B1(_00389_),
    .B2(_00390_),
    .X(_00392_));
 sky130_fd_sc_hd__a31o_1 _07012_ (.A1(net27),
    .A2(net41),
    .A3(_00277_),
    .B1(_00275_),
    .X(_00393_));
 sky130_fd_sc_hd__o21ba_1 _07013_ (.A1(_00296_),
    .A2(_00299_),
    .B1_N(_00295_),
    .X(_00394_));
 sky130_fd_sc_hd__and4_1 _07014_ (.A(net29),
    .B(net30),
    .C(net39),
    .D(net40),
    .X(_00395_));
 sky130_fd_sc_hd__a22oi_1 _07015_ (.A1(net30),
    .A2(net39),
    .B1(net40),
    .B2(net29),
    .Y(_00397_));
 sky130_fd_sc_hd__nor2_1 _07016_ (.A(_00395_),
    .B(_00397_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _07017_ (.A(net28),
    .B(net41),
    .Y(_00399_));
 sky130_fd_sc_hd__xnor2_1 _07018_ (.A(_00398_),
    .B(_00399_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand2b_1 _07019_ (.A_N(_00394_),
    .B(_00400_),
    .Y(_00401_));
 sky130_fd_sc_hd__xnor2_1 _07020_ (.A(_00394_),
    .B(_00400_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand2_1 _07021_ (.A(_00393_),
    .B(_00402_),
    .Y(_00403_));
 sky130_fd_sc_hd__xnor2_1 _07022_ (.A(_00393_),
    .B(_00402_),
    .Y(_00404_));
 sky130_fd_sc_hd__a21o_1 _07023_ (.A1(_00280_),
    .A2(_00282_),
    .B1(_00404_),
    .X(_00405_));
 sky130_fd_sc_hd__nand3_1 _07024_ (.A(_00280_),
    .B(_00282_),
    .C(_00404_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand4_2 _07025_ (.A(_00391_),
    .B(_00392_),
    .C(_00405_),
    .D(_00406_),
    .Y(_00408_));
 sky130_fd_sc_hd__a22o_1 _07026_ (.A1(_00391_),
    .A2(_00392_),
    .B1(_00405_),
    .B2(_00406_),
    .X(_00409_));
 sky130_fd_sc_hd__o211a_1 _07027_ (.A1(_00313_),
    .A2(_00315_),
    .B1(_00408_),
    .C1(_00409_),
    .X(_00410_));
 sky130_fd_sc_hd__a211oi_1 _07028_ (.A1(_00408_),
    .A2(_00409_),
    .B1(_00313_),
    .C1(_00315_),
    .Y(_00411_));
 sky130_fd_sc_hd__a211oi_1 _07029_ (.A1(_00285_),
    .A2(_00289_),
    .B1(_00410_),
    .C1(_00411_),
    .Y(_00412_));
 sky130_fd_sc_hd__o211a_1 _07030_ (.A1(_00410_),
    .A2(_00411_),
    .B1(_00285_),
    .C1(_00289_),
    .X(_00413_));
 sky130_fd_sc_hd__and4_1 _07031_ (.A(net2),
    .B(net32),
    .C(net36),
    .D(net37),
    .X(_00414_));
 sky130_fd_sc_hd__a22oi_1 _07032_ (.A1(net2),
    .A2(net36),
    .B1(net37),
    .B2(net32),
    .Y(_00415_));
 sky130_fd_sc_hd__nor2_1 _07033_ (.A(_00414_),
    .B(_00415_),
    .Y(_00416_));
 sky130_fd_sc_hd__nand2_1 _07034_ (.A(net31),
    .B(net38),
    .Y(_00417_));
 sky130_fd_sc_hd__xnor2_1 _07035_ (.A(_00416_),
    .B(_00417_),
    .Y(_00419_));
 sky130_fd_sc_hd__and4_1 _07036_ (.A(net64),
    .B(net34),
    .C(net4),
    .D(net5),
    .X(_00420_));
 sky130_fd_sc_hd__a22o_1 _07037_ (.A1(net34),
    .A2(net4),
    .B1(net5),
    .B2(net64),
    .X(_00421_));
 sky130_fd_sc_hd__and2b_1 _07038_ (.A_N(_00420_),
    .B(_00421_),
    .X(_00422_));
 sky130_fd_sc_hd__nand2_1 _07039_ (.A(net3),
    .B(net35),
    .Y(_00423_));
 sky130_fd_sc_hd__xnor2_1 _07040_ (.A(_00422_),
    .B(_00423_),
    .Y(_00424_));
 sky130_fd_sc_hd__o21ba_1 _07041_ (.A1(_00302_),
    .A2(_00304_),
    .B1_N(_00301_),
    .X(_00425_));
 sky130_fd_sc_hd__and2b_1 _07042_ (.A_N(_00425_),
    .B(_00424_),
    .X(_00426_));
 sky130_fd_sc_hd__xnor2_1 _07043_ (.A(_00424_),
    .B(_00425_),
    .Y(_00427_));
 sky130_fd_sc_hd__and2_1 _07044_ (.A(_00419_),
    .B(_00427_),
    .X(_00428_));
 sky130_fd_sc_hd__xnor2_1 _07045_ (.A(_00419_),
    .B(_00427_),
    .Y(_00430_));
 sky130_fd_sc_hd__a21o_1 _07046_ (.A1(_00325_),
    .A2(_00327_),
    .B1(_00430_),
    .X(_00431_));
 sky130_fd_sc_hd__nand3_2 _07047_ (.A(_00325_),
    .B(_00327_),
    .C(_00430_),
    .Y(_00432_));
 sky130_fd_sc_hd__o211a_1 _07048_ (.A1(_00307_),
    .A2(_00310_),
    .B1(_00431_),
    .C1(_00432_),
    .X(_00433_));
 sky130_fd_sc_hd__o211ai_2 _07049_ (.A1(_00307_),
    .A2(_00310_),
    .B1(_00431_),
    .C1(_00432_),
    .Y(_00434_));
 sky130_fd_sc_hd__a211oi_2 _07050_ (.A1(_00431_),
    .A2(_00432_),
    .B1(_00307_),
    .C1(_00310_),
    .Y(_00435_));
 sky130_fd_sc_hd__a31o_1 _07051_ (.A1(net63),
    .A2(net5),
    .A3(_00322_),
    .B1(_00319_),
    .X(_00436_));
 sky130_fd_sc_hd__o21bai_1 _07052_ (.A1(_00329_),
    .A2(_00332_),
    .B1_N(_00330_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand4_1 _07053_ (.A(net61),
    .B(net62),
    .C(net7),
    .D(net8),
    .Y(_00438_));
 sky130_fd_sc_hd__a22o_1 _07054_ (.A1(net62),
    .A2(net7),
    .B1(net8),
    .B2(net61),
    .X(_00439_));
 sky130_fd_sc_hd__nand2_1 _07055_ (.A(net63),
    .B(net6),
    .Y(_00441_));
 sky130_fd_sc_hd__nand3b_1 _07056_ (.A_N(_00441_),
    .B(_00439_),
    .C(_00438_),
    .Y(_00442_));
 sky130_fd_sc_hd__a21bo_1 _07057_ (.A1(_00438_),
    .A2(_00439_),
    .B1_N(_00441_),
    .X(_00443_));
 sky130_fd_sc_hd__and3_1 _07058_ (.A(_00437_),
    .B(_00442_),
    .C(_00443_),
    .X(_00444_));
 sky130_fd_sc_hd__a21o_1 _07059_ (.A1(_00442_),
    .A2(_00443_),
    .B1(_00437_),
    .X(_00445_));
 sky130_fd_sc_hd__and2b_1 _07060_ (.A_N(_00444_),
    .B(_00445_),
    .X(_00446_));
 sky130_fd_sc_hd__xor2_2 _07061_ (.A(_00436_),
    .B(_00446_),
    .X(_00447_));
 sky130_fd_sc_hd__nand2_1 _07062_ (.A(net60),
    .B(net9),
    .Y(_00448_));
 sky130_fd_sc_hd__and4_1 _07063_ (.A(net58),
    .B(net59),
    .C(net10),
    .D(net11),
    .X(_00449_));
 sky130_fd_sc_hd__a22oi_1 _07064_ (.A1(net59),
    .A2(net10),
    .B1(net11),
    .B2(net58),
    .Y(_00450_));
 sky130_fd_sc_hd__nor2_1 _07065_ (.A(_00449_),
    .B(_00450_),
    .Y(_00452_));
 sky130_fd_sc_hd__xnor2_1 _07066_ (.A(_00448_),
    .B(_00452_),
    .Y(_00453_));
 sky130_fd_sc_hd__nand2_1 _07067_ (.A(net55),
    .B(net13),
    .Y(_00454_));
 sky130_fd_sc_hd__and4_1 _07068_ (.A(net33),
    .B(net44),
    .C(net14),
    .D(net15),
    .X(_00455_));
 sky130_fd_sc_hd__a22oi_2 _07069_ (.A1(net44),
    .A2(net14),
    .B1(net15),
    .B2(net33),
    .Y(_00456_));
 sky130_fd_sc_hd__or3_1 _07070_ (.A(_00454_),
    .B(_00455_),
    .C(_00456_),
    .X(_00457_));
 sky130_fd_sc_hd__o21ai_1 _07071_ (.A1(_00455_),
    .A2(_00456_),
    .B1(_00454_),
    .Y(_00458_));
 sky130_fd_sc_hd__o21bai_1 _07072_ (.A1(_00335_),
    .A2(_00337_),
    .B1_N(_00336_),
    .Y(_00459_));
 sky130_fd_sc_hd__nand3_1 _07073_ (.A(_00457_),
    .B(_00458_),
    .C(_00459_),
    .Y(_00460_));
 sky130_fd_sc_hd__a21o_1 _07074_ (.A1(_00457_),
    .A2(_00458_),
    .B1(_00459_),
    .X(_00461_));
 sky130_fd_sc_hd__nand3_2 _07075_ (.A(_00453_),
    .B(_00460_),
    .C(_00461_),
    .Y(_00463_));
 sky130_fd_sc_hd__a21o_1 _07076_ (.A1(_00460_),
    .A2(_00461_),
    .B1(_00453_),
    .X(_00464_));
 sky130_fd_sc_hd__a21bo_1 _07077_ (.A1(_00334_),
    .A2(_00343_),
    .B1_N(_00341_),
    .X(_00465_));
 sky130_fd_sc_hd__nand3_4 _07078_ (.A(_00463_),
    .B(_00464_),
    .C(_00465_),
    .Y(_00466_));
 sky130_fd_sc_hd__a21o_1 _07079_ (.A1(_00463_),
    .A2(_00464_),
    .B1(_00465_),
    .X(_00467_));
 sky130_fd_sc_hd__and3_1 _07080_ (.A(_00447_),
    .B(_00466_),
    .C(_00467_),
    .X(_00468_));
 sky130_fd_sc_hd__nand3_2 _07081_ (.A(_00447_),
    .B(_00466_),
    .C(_00467_),
    .Y(_00469_));
 sky130_fd_sc_hd__a21oi_2 _07082_ (.A1(_00466_),
    .A2(_00467_),
    .B1(_00447_),
    .Y(_00470_));
 sky130_fd_sc_hd__a211oi_4 _07083_ (.A1(_00347_),
    .A2(_00350_),
    .B1(_00468_),
    .C1(_00470_),
    .Y(_00471_));
 sky130_fd_sc_hd__o211a_1 _07084_ (.A1(_00468_),
    .A2(_00470_),
    .B1(_00347_),
    .C1(_00350_),
    .X(_00472_));
 sky130_fd_sc_hd__nor4_2 _07085_ (.A(_00433_),
    .B(_00435_),
    .C(_00471_),
    .D(_00472_),
    .Y(_00474_));
 sky130_fd_sc_hd__or4_2 _07086_ (.A(_00433_),
    .B(_00435_),
    .C(_00471_),
    .D(_00472_),
    .X(_00475_));
 sky130_fd_sc_hd__o22ai_2 _07087_ (.A1(_00433_),
    .A2(_00435_),
    .B1(_00471_),
    .B2(_00472_),
    .Y(_00476_));
 sky130_fd_sc_hd__o211ai_4 _07088_ (.A1(_00352_),
    .A2(_00355_),
    .B1(_00475_),
    .C1(_00476_),
    .Y(_00477_));
 sky130_fd_sc_hd__a211o_1 _07089_ (.A1(_00475_),
    .A2(_00476_),
    .B1(_00352_),
    .C1(_00355_),
    .X(_00478_));
 sky130_fd_sc_hd__and4bb_1 _07090_ (.A_N(_00412_),
    .B_N(_00413_),
    .C(_00477_),
    .D(_00478_),
    .X(_00479_));
 sky130_fd_sc_hd__or4bb_2 _07091_ (.A(_00412_),
    .B(_00413_),
    .C_N(_00477_),
    .D_N(_00478_),
    .X(_00480_));
 sky130_fd_sc_hd__a2bb2oi_1 _07092_ (.A1_N(_00412_),
    .A2_N(_00413_),
    .B1(_00477_),
    .B2(_00478_),
    .Y(_00481_));
 sky130_fd_sc_hd__a211o_1 _07093_ (.A1(_00358_),
    .A2(_00361_),
    .B1(_00479_),
    .C1(_00481_),
    .X(_00482_));
 sky130_fd_sc_hd__o211ai_1 _07094_ (.A1(_00479_),
    .A2(_00481_),
    .B1(_00358_),
    .C1(_00361_),
    .Y(_00483_));
 sky130_fd_sc_hd__and3_1 _07095_ (.A(_00379_),
    .B(_00482_),
    .C(_00483_),
    .X(_00485_));
 sky130_fd_sc_hd__nand3_1 _07096_ (.A(_00379_),
    .B(_00482_),
    .C(_00483_),
    .Y(_00486_));
 sky130_fd_sc_hd__a21oi_1 _07097_ (.A1(_00482_),
    .A2(_00483_),
    .B1(_00379_),
    .Y(_00487_));
 sky130_fd_sc_hd__a211oi_2 _07098_ (.A1(_00363_),
    .A2(_00366_),
    .B1(_00485_),
    .C1(_00487_),
    .Y(_00488_));
 sky130_fd_sc_hd__o211a_1 _07099_ (.A1(_00485_),
    .A2(_00487_),
    .B1(_00363_),
    .C1(_00366_),
    .X(_00489_));
 sky130_fd_sc_hd__nor3_1 _07100_ (.A(_00260_),
    .B(_00488_),
    .C(_00489_),
    .Y(_00490_));
 sky130_fd_sc_hd__o21a_1 _07101_ (.A1(_00488_),
    .A2(_00489_),
    .B1(_00260_),
    .X(_00491_));
 sky130_fd_sc_hd__or2_1 _07102_ (.A(_00490_),
    .B(_00491_),
    .X(_00492_));
 sky130_fd_sc_hd__nor2_1 _07103_ (.A(_00368_),
    .B(_00492_),
    .Y(_00493_));
 sky130_fd_sc_hd__xor2_1 _07104_ (.A(_00368_),
    .B(_00492_),
    .X(_00494_));
 sky130_fd_sc_hd__and2_1 _07105_ (.A(_00371_),
    .B(_00494_),
    .X(_00496_));
 sky130_fd_sc_hd__xnor2_2 _07106_ (.A(_00371_),
    .B(_00494_),
    .Y(_00497_));
 sky130_fd_sc_hd__o21a_1 _07107_ (.A1(_00250_),
    .A2(_00252_),
    .B1(_00372_),
    .X(_00498_));
 sky130_fd_sc_hd__a21oi_1 _07108_ (.A1(_00259_),
    .A2(_00373_),
    .B1(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__xor2_1 _07109_ (.A(_00497_),
    .B(_00499_),
    .X(net79));
 sky130_fd_sc_hd__or2_1 _07110_ (.A(_00410_),
    .B(_00412_),
    .X(_00500_));
 sky130_fd_sc_hd__or2_1 _07111_ (.A(_00381_),
    .B(_00389_),
    .X(_00501_));
 sky130_fd_sc_hd__nand3_1 _07112_ (.A(_00381_),
    .B(_00389_),
    .C(_00391_),
    .Y(_00502_));
 sky130_fd_sc_hd__and2_1 _07113_ (.A(_00501_),
    .B(_00502_),
    .X(_00503_));
 sky130_fd_sc_hd__and2_1 _07114_ (.A(_00500_),
    .B(_00503_),
    .X(_00504_));
 sky130_fd_sc_hd__xnor2_1 _07115_ (.A(_00500_),
    .B(_00503_),
    .Y(_00506_));
 sky130_fd_sc_hd__and4_1 _07116_ (.A(net23),
    .B(net12),
    .C(net46),
    .D(net47),
    .X(_00507_));
 sky130_fd_sc_hd__a22o_1 _07117_ (.A1(net23),
    .A2(net46),
    .B1(net47),
    .B2(net12),
    .X(_00508_));
 sky130_fd_sc_hd__and2b_1 _07118_ (.A_N(_00507_),
    .B(_00508_),
    .X(_00509_));
 sky130_fd_sc_hd__nand2_1 _07119_ (.A(net1),
    .B(net48),
    .Y(_00510_));
 sky130_fd_sc_hd__xnor2_1 _07120_ (.A(_00509_),
    .B(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__and4_1 _07121_ (.A(net28),
    .B(net27),
    .C(net42),
    .D(net43),
    .X(_00512_));
 sky130_fd_sc_hd__a22o_1 _07122_ (.A1(net28),
    .A2(net42),
    .B1(net43),
    .B2(net27),
    .X(_00513_));
 sky130_fd_sc_hd__and2b_1 _07123_ (.A_N(_00512_),
    .B(_00513_),
    .X(_00514_));
 sky130_fd_sc_hd__nand2_1 _07124_ (.A(net26),
    .B(net45),
    .Y(_00515_));
 sky130_fd_sc_hd__xnor2_1 _07125_ (.A(_00514_),
    .B(_00515_),
    .Y(_00517_));
 sky130_fd_sc_hd__a31o_1 _07126_ (.A1(net23),
    .A2(net45),
    .A3(_00383_),
    .B1(_00382_),
    .X(_00518_));
 sky130_fd_sc_hd__and2_1 _07127_ (.A(_00517_),
    .B(_00518_),
    .X(_00519_));
 sky130_fd_sc_hd__xor2_1 _07128_ (.A(_00517_),
    .B(_00518_),
    .X(_00520_));
 sky130_fd_sc_hd__and2_1 _07129_ (.A(_00511_),
    .B(_00520_),
    .X(_00521_));
 sky130_fd_sc_hd__nor2_1 _07130_ (.A(_00511_),
    .B(_00520_),
    .Y(_00522_));
 sky130_fd_sc_hd__or2_1 _07131_ (.A(_00521_),
    .B(_00522_),
    .X(_00523_));
 sky130_fd_sc_hd__a31o_1 _07132_ (.A1(net28),
    .A2(net41),
    .A3(_00398_),
    .B1(_00395_),
    .X(_00524_));
 sky130_fd_sc_hd__o21bai_1 _07133_ (.A1(_00415_),
    .A2(_00417_),
    .B1_N(_00414_),
    .Y(_00525_));
 sky130_fd_sc_hd__nand4_1 _07134_ (.A(net30),
    .B(net31),
    .C(net39),
    .D(net40),
    .Y(_00526_));
 sky130_fd_sc_hd__a22o_1 _07135_ (.A1(net31),
    .A2(net39),
    .B1(net40),
    .B2(net30),
    .X(_00528_));
 sky130_fd_sc_hd__nand2_1 _07136_ (.A(net29),
    .B(net41),
    .Y(_00529_));
 sky130_fd_sc_hd__nand3b_1 _07137_ (.A_N(_00529_),
    .B(_00528_),
    .C(_00526_),
    .Y(_00530_));
 sky130_fd_sc_hd__a21bo_1 _07138_ (.A1(_00526_),
    .A2(_00528_),
    .B1_N(_00529_),
    .X(_00531_));
 sky130_fd_sc_hd__and3_1 _07139_ (.A(_00525_),
    .B(_00530_),
    .C(_00531_),
    .X(_00532_));
 sky130_fd_sc_hd__a21o_1 _07140_ (.A1(_00530_),
    .A2(_00531_),
    .B1(_00525_),
    .X(_00533_));
 sky130_fd_sc_hd__and2b_1 _07141_ (.A_N(_00532_),
    .B(_00533_),
    .X(_00534_));
 sky130_fd_sc_hd__xnor2_1 _07142_ (.A(_00524_),
    .B(_00534_),
    .Y(_00535_));
 sky130_fd_sc_hd__a21oi_2 _07143_ (.A1(_00401_),
    .A2(_00403_),
    .B1(_00535_),
    .Y(_00536_));
 sky130_fd_sc_hd__inv_2 _07144_ (.A(_00536_),
    .Y(_00537_));
 sky130_fd_sc_hd__and3_1 _07145_ (.A(_00401_),
    .B(_00403_),
    .C(_00535_),
    .X(_00539_));
 sky130_fd_sc_hd__nor3_1 _07146_ (.A(_00523_),
    .B(_00536_),
    .C(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__or3_1 _07147_ (.A(_00523_),
    .B(_00536_),
    .C(_00539_),
    .X(_00541_));
 sky130_fd_sc_hd__o21a_1 _07148_ (.A1(_00536_),
    .A2(_00539_),
    .B1(_00523_),
    .X(_00542_));
 sky130_fd_sc_hd__a211oi_2 _07149_ (.A1(_00431_),
    .A2(_00434_),
    .B1(_00540_),
    .C1(_00542_),
    .Y(_00543_));
 sky130_fd_sc_hd__o211a_1 _07150_ (.A1(_00540_),
    .A2(_00542_),
    .B1(_00431_),
    .C1(_00434_),
    .X(_00544_));
 sky130_fd_sc_hd__a211oi_2 _07151_ (.A1(_00405_),
    .A2(_00408_),
    .B1(_00543_),
    .C1(_00544_),
    .Y(_00545_));
 sky130_fd_sc_hd__o211a_1 _07152_ (.A1(_00543_),
    .A2(_00544_),
    .B1(_00405_),
    .C1(_00408_),
    .X(_00546_));
 sky130_fd_sc_hd__a21o_1 _07153_ (.A1(_00436_),
    .A2(_00445_),
    .B1(_00444_),
    .X(_00547_));
 sky130_fd_sc_hd__and4_1 _07154_ (.A(net2),
    .B(net3),
    .C(net36),
    .D(net37),
    .X(_00548_));
 sky130_fd_sc_hd__a22o_1 _07155_ (.A1(net3),
    .A2(net36),
    .B1(net37),
    .B2(net2),
    .X(_00550_));
 sky130_fd_sc_hd__and2b_1 _07156_ (.A_N(_00548_),
    .B(_00550_),
    .X(_00551_));
 sky130_fd_sc_hd__nand2_1 _07157_ (.A(net32),
    .B(net38),
    .Y(_00552_));
 sky130_fd_sc_hd__xnor2_1 _07158_ (.A(_00551_),
    .B(_00552_),
    .Y(_00553_));
 sky130_fd_sc_hd__and4_1 _07159_ (.A(net64),
    .B(net34),
    .C(net5),
    .D(net6),
    .X(_00554_));
 sky130_fd_sc_hd__a22oi_2 _07160_ (.A1(net34),
    .A2(net5),
    .B1(net6),
    .B2(net64),
    .Y(_00555_));
 sky130_fd_sc_hd__nand2_1 _07161_ (.A(net35),
    .B(net4),
    .Y(_00556_));
 sky130_fd_sc_hd__or3_1 _07162_ (.A(_00554_),
    .B(_00555_),
    .C(_00556_),
    .X(_00557_));
 sky130_fd_sc_hd__o21ai_1 _07163_ (.A1(_00554_),
    .A2(_00555_),
    .B1(_00556_),
    .Y(_00558_));
 sky130_fd_sc_hd__a31o_1 _07164_ (.A1(net3),
    .A2(net35),
    .A3(_00421_),
    .B1(_00420_),
    .X(_00559_));
 sky130_fd_sc_hd__nand3_2 _07165_ (.A(_00557_),
    .B(_00558_),
    .C(_00559_),
    .Y(_00561_));
 sky130_fd_sc_hd__a21o_1 _07166_ (.A1(_00557_),
    .A2(_00558_),
    .B1(_00559_),
    .X(_00562_));
 sky130_fd_sc_hd__nand3_2 _07167_ (.A(_00553_),
    .B(_00561_),
    .C(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__a21o_1 _07168_ (.A1(_00561_),
    .A2(_00562_),
    .B1(_00553_),
    .X(_00564_));
 sky130_fd_sc_hd__nand3_2 _07169_ (.A(_00547_),
    .B(_00563_),
    .C(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__a21o_1 _07170_ (.A1(_00563_),
    .A2(_00564_),
    .B1(_00547_),
    .X(_00566_));
 sky130_fd_sc_hd__o211ai_2 _07171_ (.A1(_00426_),
    .A2(_00428_),
    .B1(_00565_),
    .C1(_00566_),
    .Y(_00567_));
 sky130_fd_sc_hd__a211o_1 _07172_ (.A1(_00565_),
    .A2(_00566_),
    .B1(_00426_),
    .C1(_00428_),
    .X(_00568_));
 sky130_fd_sc_hd__nand2_1 _07173_ (.A(_00567_),
    .B(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_1 _07174_ (.A(_00438_),
    .B(_00442_),
    .Y(_00570_));
 sky130_fd_sc_hd__o21bai_1 _07175_ (.A1(_00448_),
    .A2(_00450_),
    .B1_N(_00449_),
    .Y(_00572_));
 sky130_fd_sc_hd__and4_1 _07176_ (.A(net61),
    .B(net62),
    .C(net8),
    .D(net9),
    .X(_00573_));
 sky130_fd_sc_hd__a22oi_1 _07177_ (.A1(net62),
    .A2(net8),
    .B1(net9),
    .B2(net61),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _07178_ (.A(net63),
    .B(net7),
    .Y(_00575_));
 sky130_fd_sc_hd__or3_1 _07179_ (.A(_00573_),
    .B(_00574_),
    .C(_00575_),
    .X(_00576_));
 sky130_fd_sc_hd__o21ai_1 _07180_ (.A1(_00573_),
    .A2(_00574_),
    .B1(_00575_),
    .Y(_00577_));
 sky130_fd_sc_hd__and3_1 _07181_ (.A(_00572_),
    .B(_00576_),
    .C(_00577_),
    .X(_00578_));
 sky130_fd_sc_hd__a21o_1 _07182_ (.A1(_00576_),
    .A2(_00577_),
    .B1(_00572_),
    .X(_00579_));
 sky130_fd_sc_hd__and2b_1 _07183_ (.A_N(_00578_),
    .B(_00579_),
    .X(_00580_));
 sky130_fd_sc_hd__xor2_1 _07184_ (.A(_00570_),
    .B(_00580_),
    .X(_00581_));
 sky130_fd_sc_hd__nand2_1 _07185_ (.A(net60),
    .B(net10),
    .Y(_00583_));
 sky130_fd_sc_hd__and4_1 _07186_ (.A(net58),
    .B(net59),
    .C(net11),
    .D(net13),
    .X(_00584_));
 sky130_fd_sc_hd__a22oi_1 _07187_ (.A1(net59),
    .A2(net11),
    .B1(net13),
    .B2(net58),
    .Y(_00585_));
 sky130_fd_sc_hd__nor2_1 _07188_ (.A(_00584_),
    .B(_00585_),
    .Y(_00586_));
 sky130_fd_sc_hd__xnor2_1 _07189_ (.A(_00583_),
    .B(_00586_),
    .Y(_00587_));
 sky130_fd_sc_hd__nand2_1 _07190_ (.A(net55),
    .B(net14),
    .Y(_00588_));
 sky130_fd_sc_hd__and4_1 _07191_ (.A(net33),
    .B(net44),
    .C(net15),
    .D(net16),
    .X(_00589_));
 sky130_fd_sc_hd__a22oi_2 _07192_ (.A1(net44),
    .A2(net15),
    .B1(net16),
    .B2(net33),
    .Y(_00590_));
 sky130_fd_sc_hd__or3_1 _07193_ (.A(_00588_),
    .B(_00589_),
    .C(_00590_),
    .X(_00591_));
 sky130_fd_sc_hd__o21ai_1 _07194_ (.A1(_00589_),
    .A2(_00590_),
    .B1(_00588_),
    .Y(_00592_));
 sky130_fd_sc_hd__o21bai_1 _07195_ (.A1(_00454_),
    .A2(_00456_),
    .B1_N(_00455_),
    .Y(_00594_));
 sky130_fd_sc_hd__nand3_1 _07196_ (.A(_00591_),
    .B(_00592_),
    .C(_00594_),
    .Y(_00595_));
 sky130_fd_sc_hd__a21o_1 _07197_ (.A1(_00591_),
    .A2(_00592_),
    .B1(_00594_),
    .X(_00596_));
 sky130_fd_sc_hd__nand3_1 _07198_ (.A(_00587_),
    .B(_00595_),
    .C(_00596_),
    .Y(_00597_));
 sky130_fd_sc_hd__a21o_1 _07199_ (.A1(_00595_),
    .A2(_00596_),
    .B1(_00587_),
    .X(_00598_));
 sky130_fd_sc_hd__a21bo_1 _07200_ (.A1(_00453_),
    .A2(_00461_),
    .B1_N(_00460_),
    .X(_00599_));
 sky130_fd_sc_hd__nand3_2 _07201_ (.A(_00597_),
    .B(_00598_),
    .C(_00599_),
    .Y(_00600_));
 sky130_fd_sc_hd__a21o_1 _07202_ (.A1(_00597_),
    .A2(_00598_),
    .B1(_00599_),
    .X(_00601_));
 sky130_fd_sc_hd__and3_1 _07203_ (.A(_00581_),
    .B(_00600_),
    .C(_00601_),
    .X(_00602_));
 sky130_fd_sc_hd__nand3_1 _07204_ (.A(_00581_),
    .B(_00600_),
    .C(_00601_),
    .Y(_00603_));
 sky130_fd_sc_hd__a21oi_2 _07205_ (.A1(_00600_),
    .A2(_00601_),
    .B1(_00581_),
    .Y(_00605_));
 sky130_fd_sc_hd__a211oi_4 _07206_ (.A1(_00466_),
    .A2(_00469_),
    .B1(_00602_),
    .C1(_00605_),
    .Y(_00606_));
 sky130_fd_sc_hd__o211a_1 _07207_ (.A1(_00602_),
    .A2(_00605_),
    .B1(_00466_),
    .C1(_00469_),
    .X(_00607_));
 sky130_fd_sc_hd__nor3_1 _07208_ (.A(_00569_),
    .B(_00606_),
    .C(_00607_),
    .Y(_00608_));
 sky130_fd_sc_hd__or3_2 _07209_ (.A(_00569_),
    .B(_00606_),
    .C(_00607_),
    .X(_00609_));
 sky130_fd_sc_hd__o21ai_2 _07210_ (.A1(_00606_),
    .A2(_00607_),
    .B1(_00569_),
    .Y(_00610_));
 sky130_fd_sc_hd__o211ai_4 _07211_ (.A1(_00471_),
    .A2(_00474_),
    .B1(_00609_),
    .C1(_00610_),
    .Y(_00611_));
 sky130_fd_sc_hd__a211o_1 _07212_ (.A1(_00609_),
    .A2(_00610_),
    .B1(_00471_),
    .C1(_00474_),
    .X(_00612_));
 sky130_fd_sc_hd__and4bb_1 _07213_ (.A_N(_00545_),
    .B_N(_00546_),
    .C(_00611_),
    .D(_00612_),
    .X(_00613_));
 sky130_fd_sc_hd__or4bb_1 _07214_ (.A(_00545_),
    .B(_00546_),
    .C_N(_00611_),
    .D_N(_00612_),
    .X(_00614_));
 sky130_fd_sc_hd__a2bb2oi_2 _07215_ (.A1_N(_00545_),
    .A2_N(_00546_),
    .B1(_00611_),
    .B2(_00612_),
    .Y(_00616_));
 sky130_fd_sc_hd__a211oi_4 _07216_ (.A1(_00477_),
    .A2(_00480_),
    .B1(_00613_),
    .C1(_00616_),
    .Y(_00617_));
 sky130_fd_sc_hd__o211a_1 _07217_ (.A1(_00613_),
    .A2(_00616_),
    .B1(_00477_),
    .C1(_00480_),
    .X(_00618_));
 sky130_fd_sc_hd__nor3_2 _07218_ (.A(_00506_),
    .B(_00617_),
    .C(_00618_),
    .Y(_00619_));
 sky130_fd_sc_hd__o21a_1 _07219_ (.A1(_00617_),
    .A2(_00618_),
    .B1(_00506_),
    .X(_00620_));
 sky130_fd_sc_hd__a211oi_1 _07220_ (.A1(_00482_),
    .A2(_00486_),
    .B1(_00619_),
    .C1(_00620_),
    .Y(_00621_));
 sky130_fd_sc_hd__a211o_1 _07221_ (.A1(_00482_),
    .A2(_00486_),
    .B1(_00619_),
    .C1(_00620_),
    .X(_00622_));
 sky130_fd_sc_hd__o211ai_1 _07222_ (.A1(_00619_),
    .A2(_00620_),
    .B1(_00482_),
    .C1(_00486_),
    .Y(_00623_));
 sky130_fd_sc_hd__and3_1 _07223_ (.A(_00377_),
    .B(_00622_),
    .C(_00623_),
    .X(_00624_));
 sky130_fd_sc_hd__nand3_1 _07224_ (.A(_00377_),
    .B(_00622_),
    .C(_00623_),
    .Y(_00625_));
 sky130_fd_sc_hd__a21o_1 _07225_ (.A1(_00622_),
    .A2(_00623_),
    .B1(_00377_),
    .X(_00627_));
 sky130_fd_sc_hd__o211a_1 _07226_ (.A1(_00488_),
    .A2(_00490_),
    .B1(_00625_),
    .C1(_00627_),
    .X(_00628_));
 sky130_fd_sc_hd__a211oi_1 _07227_ (.A1(_00625_),
    .A2(_00627_),
    .B1(_00488_),
    .C1(_00490_),
    .Y(_00629_));
 sky130_fd_sc_hd__nor2_1 _07228_ (.A(_00628_),
    .B(_00629_),
    .Y(_00630_));
 sky130_fd_sc_hd__xor2_1 _07229_ (.A(_00493_),
    .B(_00630_),
    .X(_00631_));
 sky130_fd_sc_hd__o21ba_1 _07230_ (.A1(_00497_),
    .A2(_00499_),
    .B1_N(_00496_),
    .X(_00632_));
 sky130_fd_sc_hd__xnor2_1 _07231_ (.A(_00631_),
    .B(_00632_),
    .Y(net80));
 sky130_fd_sc_hd__or2_1 _07232_ (.A(_00543_),
    .B(_00545_),
    .X(_00633_));
 sky130_fd_sc_hd__a31o_1 _07233_ (.A1(net1),
    .A2(net48),
    .A3(_00508_),
    .B1(_00507_),
    .X(_00634_));
 sky130_fd_sc_hd__and3_1 _07234_ (.A(net1),
    .B(net49),
    .C(_00634_),
    .X(_00635_));
 sky130_fd_sc_hd__a21oi_1 _07235_ (.A1(net1),
    .A2(net49),
    .B1(_00634_),
    .Y(_00637_));
 sky130_fd_sc_hd__nor2_1 _07236_ (.A(_00635_),
    .B(_00637_),
    .Y(_00638_));
 sky130_fd_sc_hd__o21ai_1 _07237_ (.A1(_00519_),
    .A2(_00521_),
    .B1(_00638_),
    .Y(_00639_));
 sky130_fd_sc_hd__or3_1 _07238_ (.A(_00519_),
    .B(_00521_),
    .C(_00638_),
    .X(_00640_));
 sky130_fd_sc_hd__and2_1 _07239_ (.A(_00639_),
    .B(_00640_),
    .X(_00641_));
 sky130_fd_sc_hd__and2b_1 _07240_ (.A_N(_00501_),
    .B(_00641_),
    .X(_00642_));
 sky130_fd_sc_hd__xnor2_1 _07241_ (.A(_00501_),
    .B(_00641_),
    .Y(_00643_));
 sky130_fd_sc_hd__nand2_1 _07242_ (.A(_00633_),
    .B(_00643_),
    .Y(_00644_));
 sky130_fd_sc_hd__xnor2_1 _07243_ (.A(_00633_),
    .B(_00643_),
    .Y(_00645_));
 sky130_fd_sc_hd__and4_1 _07244_ (.A(net26),
    .B(net23),
    .C(net46),
    .D(net47),
    .X(_00646_));
 sky130_fd_sc_hd__a22oi_1 _07245_ (.A1(net26),
    .A2(net46),
    .B1(net47),
    .B2(net23),
    .Y(_00648_));
 sky130_fd_sc_hd__nor2_1 _07246_ (.A(_00646_),
    .B(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__nand2_1 _07247_ (.A(net12),
    .B(net48),
    .Y(_00650_));
 sky130_fd_sc_hd__xnor2_1 _07248_ (.A(_00649_),
    .B(_00650_),
    .Y(_00651_));
 sky130_fd_sc_hd__and4_1 _07249_ (.A(net28),
    .B(net29),
    .C(net42),
    .D(net43),
    .X(_00652_));
 sky130_fd_sc_hd__a22oi_2 _07250_ (.A1(net29),
    .A2(net42),
    .B1(net43),
    .B2(net28),
    .Y(_00653_));
 sky130_fd_sc_hd__nand2_1 _07251_ (.A(net27),
    .B(net45),
    .Y(_00654_));
 sky130_fd_sc_hd__or3_1 _07252_ (.A(_00652_),
    .B(_00653_),
    .C(_00654_),
    .X(_00655_));
 sky130_fd_sc_hd__o21ai_1 _07253_ (.A1(_00652_),
    .A2(_00653_),
    .B1(_00654_),
    .Y(_00656_));
 sky130_fd_sc_hd__a31o_1 _07254_ (.A1(net26),
    .A2(net45),
    .A3(_00513_),
    .B1(_00512_),
    .X(_00657_));
 sky130_fd_sc_hd__and3_1 _07255_ (.A(_00655_),
    .B(_00656_),
    .C(_00657_),
    .X(_00659_));
 sky130_fd_sc_hd__a21oi_1 _07256_ (.A1(_00655_),
    .A2(_00656_),
    .B1(_00657_),
    .Y(_00660_));
 sky130_fd_sc_hd__nor3b_1 _07257_ (.A(_00659_),
    .B(_00660_),
    .C_N(_00651_),
    .Y(_00661_));
 sky130_fd_sc_hd__o21ba_1 _07258_ (.A1(_00659_),
    .A2(_00660_),
    .B1_N(_00651_),
    .X(_00662_));
 sky130_fd_sc_hd__or2_1 _07259_ (.A(_00661_),
    .B(_00662_),
    .X(_00663_));
 sky130_fd_sc_hd__nand2_1 _07260_ (.A(_00526_),
    .B(_00530_),
    .Y(_00664_));
 sky130_fd_sc_hd__a31o_1 _07261_ (.A1(net32),
    .A2(net38),
    .A3(_00550_),
    .B1(_00548_),
    .X(_00665_));
 sky130_fd_sc_hd__nand4_1 _07262_ (.A(net31),
    .B(net32),
    .C(net39),
    .D(net40),
    .Y(_00666_));
 sky130_fd_sc_hd__a22o_1 _07263_ (.A1(net32),
    .A2(net39),
    .B1(net40),
    .B2(net31),
    .X(_00667_));
 sky130_fd_sc_hd__nand2_1 _07264_ (.A(net30),
    .B(net41),
    .Y(_00668_));
 sky130_fd_sc_hd__nand3b_1 _07265_ (.A_N(_00668_),
    .B(_00667_),
    .C(_00666_),
    .Y(_00670_));
 sky130_fd_sc_hd__a21bo_1 _07266_ (.A1(_00666_),
    .A2(_00667_),
    .B1_N(_00668_),
    .X(_00671_));
 sky130_fd_sc_hd__nand3_1 _07267_ (.A(_00665_),
    .B(_00670_),
    .C(_00671_),
    .Y(_00672_));
 sky130_fd_sc_hd__a21o_1 _07268_ (.A1(_00670_),
    .A2(_00671_),
    .B1(_00665_),
    .X(_00673_));
 sky130_fd_sc_hd__nand3_1 _07269_ (.A(_00664_),
    .B(_00672_),
    .C(_00673_),
    .Y(_00674_));
 sky130_fd_sc_hd__a21o_1 _07270_ (.A1(_00672_),
    .A2(_00673_),
    .B1(_00664_),
    .X(_00675_));
 sky130_fd_sc_hd__a21o_1 _07271_ (.A1(_00524_),
    .A2(_00533_),
    .B1(_00532_),
    .X(_00676_));
 sky130_fd_sc_hd__and3_1 _07272_ (.A(_00674_),
    .B(_00675_),
    .C(_00676_),
    .X(_00677_));
 sky130_fd_sc_hd__inv_2 _07273_ (.A(_00677_),
    .Y(_00678_));
 sky130_fd_sc_hd__a21oi_1 _07274_ (.A1(_00674_),
    .A2(_00675_),
    .B1(_00676_),
    .Y(_00679_));
 sky130_fd_sc_hd__nor3_1 _07275_ (.A(_00663_),
    .B(_00677_),
    .C(_00679_),
    .Y(_00681_));
 sky130_fd_sc_hd__or3_1 _07276_ (.A(_00663_),
    .B(_00677_),
    .C(_00679_),
    .X(_00682_));
 sky130_fd_sc_hd__o21a_1 _07277_ (.A1(_00677_),
    .A2(_00679_),
    .B1(_00663_),
    .X(_00683_));
 sky130_fd_sc_hd__a211oi_2 _07278_ (.A1(_00565_),
    .A2(_00567_),
    .B1(_00681_),
    .C1(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__o211a_1 _07279_ (.A1(_00681_),
    .A2(_00683_),
    .B1(_00565_),
    .C1(_00567_),
    .X(_00685_));
 sky130_fd_sc_hd__a211oi_2 _07280_ (.A1(_00537_),
    .A2(_00541_),
    .B1(_00684_),
    .C1(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__o211a_1 _07281_ (.A1(_00684_),
    .A2(_00685_),
    .B1(_00537_),
    .C1(_00541_),
    .X(_00687_));
 sky130_fd_sc_hd__a21o_1 _07282_ (.A1(_00570_),
    .A2(_00579_),
    .B1(_00578_),
    .X(_00688_));
 sky130_fd_sc_hd__and4_1 _07283_ (.A(net3),
    .B(net4),
    .C(net36),
    .D(net37),
    .X(_00689_));
 sky130_fd_sc_hd__a22o_1 _07284_ (.A1(net4),
    .A2(net36),
    .B1(net37),
    .B2(net3),
    .X(_00690_));
 sky130_fd_sc_hd__and2b_1 _07285_ (.A_N(_00689_),
    .B(_00690_),
    .X(_00692_));
 sky130_fd_sc_hd__nand2_1 _07286_ (.A(net2),
    .B(net38),
    .Y(_00693_));
 sky130_fd_sc_hd__xnor2_1 _07287_ (.A(_00692_),
    .B(_00693_),
    .Y(_00694_));
 sky130_fd_sc_hd__nand4_1 _07288_ (.A(net64),
    .B(net34),
    .C(net6),
    .D(net7),
    .Y(_00695_));
 sky130_fd_sc_hd__a22o_1 _07289_ (.A1(net34),
    .A2(net6),
    .B1(net7),
    .B2(net64),
    .X(_00696_));
 sky130_fd_sc_hd__nand2_1 _07290_ (.A(net35),
    .B(net5),
    .Y(_00697_));
 sky130_fd_sc_hd__nand3b_1 _07291_ (.A_N(_00697_),
    .B(_00696_),
    .C(_00695_),
    .Y(_00698_));
 sky130_fd_sc_hd__a21bo_1 _07292_ (.A1(_00695_),
    .A2(_00696_),
    .B1_N(_00697_),
    .X(_00699_));
 sky130_fd_sc_hd__o21bai_1 _07293_ (.A1(_00555_),
    .A2(_00556_),
    .B1_N(_00554_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand3_2 _07294_ (.A(_00698_),
    .B(_00699_),
    .C(_00700_),
    .Y(_00701_));
 sky130_fd_sc_hd__a21o_1 _07295_ (.A1(_00698_),
    .A2(_00699_),
    .B1(_00700_),
    .X(_00703_));
 sky130_fd_sc_hd__nand3_2 _07296_ (.A(_00694_),
    .B(_00701_),
    .C(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__a21o_1 _07297_ (.A1(_00701_),
    .A2(_00703_),
    .B1(_00694_),
    .X(_00705_));
 sky130_fd_sc_hd__and3_1 _07298_ (.A(_00688_),
    .B(_00704_),
    .C(_00705_),
    .X(_00706_));
 sky130_fd_sc_hd__a21oi_1 _07299_ (.A1(_00704_),
    .A2(_00705_),
    .B1(_00688_),
    .Y(_00707_));
 sky130_fd_sc_hd__a211oi_2 _07300_ (.A1(_00561_),
    .A2(_00563_),
    .B1(_00706_),
    .C1(_00707_),
    .Y(_00708_));
 sky130_fd_sc_hd__o211a_1 _07301_ (.A1(_00706_),
    .A2(_00707_),
    .B1(_00561_),
    .C1(_00563_),
    .X(_00709_));
 sky130_fd_sc_hd__and2b_1 _07302_ (.A_N(_00573_),
    .B(_00576_),
    .X(_00710_));
 sky130_fd_sc_hd__o21ba_1 _07303_ (.A1(_00583_),
    .A2(_00585_),
    .B1_N(_00584_),
    .X(_00711_));
 sky130_fd_sc_hd__and4_1 _07304_ (.A(net61),
    .B(net62),
    .C(net9),
    .D(net10),
    .X(_00712_));
 sky130_fd_sc_hd__a22oi_1 _07305_ (.A1(net62),
    .A2(net9),
    .B1(net10),
    .B2(net61),
    .Y(_00714_));
 sky130_fd_sc_hd__nor2_1 _07306_ (.A(_00712_),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__nand2_1 _07307_ (.A(net63),
    .B(net8),
    .Y(_00716_));
 sky130_fd_sc_hd__xnor2_1 _07308_ (.A(_00715_),
    .B(_00716_),
    .Y(_00717_));
 sky130_fd_sc_hd__nand2b_1 _07309_ (.A_N(_00711_),
    .B(_00717_),
    .Y(_00718_));
 sky130_fd_sc_hd__xnor2_1 _07310_ (.A(_00711_),
    .B(_00717_),
    .Y(_00719_));
 sky130_fd_sc_hd__nand2b_1 _07311_ (.A_N(_00710_),
    .B(_00719_),
    .Y(_00720_));
 sky130_fd_sc_hd__xnor2_1 _07312_ (.A(_00710_),
    .B(_00719_),
    .Y(_00721_));
 sky130_fd_sc_hd__and4_1 _07313_ (.A(net58),
    .B(net59),
    .C(net13),
    .D(net14),
    .X(_00722_));
 sky130_fd_sc_hd__a22oi_1 _07314_ (.A1(net59),
    .A2(net13),
    .B1(net14),
    .B2(net58),
    .Y(_00723_));
 sky130_fd_sc_hd__nor2_1 _07315_ (.A(_00722_),
    .B(_00723_),
    .Y(_00725_));
 sky130_fd_sc_hd__nand2_1 _07316_ (.A(net60),
    .B(net11),
    .Y(_00726_));
 sky130_fd_sc_hd__xnor2_1 _07317_ (.A(_00725_),
    .B(_00726_),
    .Y(_00727_));
 sky130_fd_sc_hd__nand2_1 _07318_ (.A(net55),
    .B(net15),
    .Y(_00728_));
 sky130_fd_sc_hd__and4_1 _07319_ (.A(net33),
    .B(net44),
    .C(net16),
    .D(net17),
    .X(_00729_));
 sky130_fd_sc_hd__a22oi_2 _07320_ (.A1(net44),
    .A2(net16),
    .B1(net17),
    .B2(net33),
    .Y(_00730_));
 sky130_fd_sc_hd__or3_1 _07321_ (.A(_00728_),
    .B(_00729_),
    .C(_00730_),
    .X(_00731_));
 sky130_fd_sc_hd__o21ai_1 _07322_ (.A1(_00729_),
    .A2(_00730_),
    .B1(_00728_),
    .Y(_00732_));
 sky130_fd_sc_hd__o21bai_1 _07323_ (.A1(_00588_),
    .A2(_00590_),
    .B1_N(_00589_),
    .Y(_00733_));
 sky130_fd_sc_hd__nand3_1 _07324_ (.A(_00731_),
    .B(_00732_),
    .C(_00733_),
    .Y(_00734_));
 sky130_fd_sc_hd__a21o_1 _07325_ (.A1(_00731_),
    .A2(_00732_),
    .B1(_00733_),
    .X(_00736_));
 sky130_fd_sc_hd__nand3_1 _07326_ (.A(_00727_),
    .B(_00734_),
    .C(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__a21o_1 _07327_ (.A1(_00734_),
    .A2(_00736_),
    .B1(_00727_),
    .X(_00738_));
 sky130_fd_sc_hd__a21bo_1 _07328_ (.A1(_00587_),
    .A2(_00596_),
    .B1_N(_00595_),
    .X(_00739_));
 sky130_fd_sc_hd__nand3_4 _07329_ (.A(_00737_),
    .B(_00738_),
    .C(_00739_),
    .Y(_00740_));
 sky130_fd_sc_hd__a21o_1 _07330_ (.A1(_00737_),
    .A2(_00738_),
    .B1(_00739_),
    .X(_00741_));
 sky130_fd_sc_hd__and3_1 _07331_ (.A(_00721_),
    .B(_00740_),
    .C(_00741_),
    .X(_00742_));
 sky130_fd_sc_hd__nand3_2 _07332_ (.A(_00721_),
    .B(_00740_),
    .C(_00741_),
    .Y(_00743_));
 sky130_fd_sc_hd__a21oi_1 _07333_ (.A1(_00740_),
    .A2(_00741_),
    .B1(_00721_),
    .Y(_00744_));
 sky130_fd_sc_hd__a211o_1 _07334_ (.A1(_00600_),
    .A2(_00603_),
    .B1(_00742_),
    .C1(_00744_),
    .X(_00745_));
 sky130_fd_sc_hd__o211ai_1 _07335_ (.A1(_00742_),
    .A2(_00744_),
    .B1(_00600_),
    .C1(_00603_),
    .Y(_00747_));
 sky130_fd_sc_hd__or4bb_2 _07336_ (.A(_00708_),
    .B(_00709_),
    .C_N(_00745_),
    .D_N(_00747_),
    .X(_00748_));
 sky130_fd_sc_hd__a2bb2o_1 _07337_ (.A1_N(_00708_),
    .A2_N(_00709_),
    .B1(_00745_),
    .B2(_00747_),
    .X(_00749_));
 sky130_fd_sc_hd__o211a_1 _07338_ (.A1(_00606_),
    .A2(_00608_),
    .B1(_00748_),
    .C1(_00749_),
    .X(_00750_));
 sky130_fd_sc_hd__a211oi_2 _07339_ (.A1(_00748_),
    .A2(_00749_),
    .B1(_00606_),
    .C1(_00608_),
    .Y(_00751_));
 sky130_fd_sc_hd__nor4_2 _07340_ (.A(_00686_),
    .B(_00687_),
    .C(_00750_),
    .D(_00751_),
    .Y(_00752_));
 sky130_fd_sc_hd__o22a_1 _07341_ (.A1(_00686_),
    .A2(_00687_),
    .B1(_00750_),
    .B2(_00751_),
    .X(_00753_));
 sky130_fd_sc_hd__a211oi_2 _07342_ (.A1(_00611_),
    .A2(_00614_),
    .B1(_00752_),
    .C1(_00753_),
    .Y(_00754_));
 sky130_fd_sc_hd__o211a_1 _07343_ (.A1(_00752_),
    .A2(_00753_),
    .B1(_00611_),
    .C1(_00614_),
    .X(_00755_));
 sky130_fd_sc_hd__nor3_1 _07344_ (.A(_00645_),
    .B(_00754_),
    .C(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__or3_1 _07345_ (.A(_00645_),
    .B(_00754_),
    .C(_00755_),
    .X(_00758_));
 sky130_fd_sc_hd__o21ai_1 _07346_ (.A1(_00754_),
    .A2(_00755_),
    .B1(_00645_),
    .Y(_00759_));
 sky130_fd_sc_hd__o211a_1 _07347_ (.A1(_00617_),
    .A2(_00619_),
    .B1(_00758_),
    .C1(_00759_),
    .X(_00760_));
 sky130_fd_sc_hd__o211ai_1 _07348_ (.A1(_00617_),
    .A2(_00619_),
    .B1(_00758_),
    .C1(_00759_),
    .Y(_00761_));
 sky130_fd_sc_hd__a211o_1 _07349_ (.A1(_00758_),
    .A2(_00759_),
    .B1(_00617_),
    .C1(_00619_),
    .X(_00762_));
 sky130_fd_sc_hd__and3_1 _07350_ (.A(_00504_),
    .B(_00761_),
    .C(_00762_),
    .X(_00763_));
 sky130_fd_sc_hd__nand3_1 _07351_ (.A(_00504_),
    .B(_00761_),
    .C(_00762_),
    .Y(_00764_));
 sky130_fd_sc_hd__a21o_1 _07352_ (.A1(_00761_),
    .A2(_00762_),
    .B1(_00504_),
    .X(_00765_));
 sky130_fd_sc_hd__o211a_1 _07353_ (.A1(_00621_),
    .A2(_00624_),
    .B1(_00764_),
    .C1(_00765_),
    .X(_00766_));
 sky130_fd_sc_hd__a211o_1 _07354_ (.A1(_00764_),
    .A2(_00765_),
    .B1(_00621_),
    .C1(_00624_),
    .X(_00767_));
 sky130_fd_sc_hd__and2b_1 _07355_ (.A_N(_00766_),
    .B(_00767_),
    .X(_00769_));
 sky130_fd_sc_hd__and3b_1 _07356_ (.A_N(_00766_),
    .B(_00767_),
    .C(_00628_),
    .X(_00770_));
 sky130_fd_sc_hd__xnor2_1 _07357_ (.A(_00628_),
    .B(_00769_),
    .Y(_00771_));
 sky130_fd_sc_hd__and4bb_1 _07358_ (.A_N(_00254_),
    .B_N(_00497_),
    .C(_00631_),
    .D(_00373_),
    .X(_00772_));
 sky130_fd_sc_hd__o21a_1 _07359_ (.A1(_00493_),
    .A2(_00496_),
    .B1(_00630_),
    .X(_00773_));
 sky130_fd_sc_hd__and3b_1 _07360_ (.A_N(_00497_),
    .B(_00498_),
    .C(_00631_),
    .X(_00774_));
 sky130_fd_sc_hd__a211o_1 _07361_ (.A1(_00257_),
    .A2(_00772_),
    .B1(_00773_),
    .C1(_00774_),
    .X(_00775_));
 sky130_fd_sc_hd__and3_1 _07362_ (.A(_00047_),
    .B(_00255_),
    .C(_00772_),
    .X(_00776_));
 sky130_fd_sc_hd__a21oi_2 _07363_ (.A1(_05524_),
    .A2(_00776_),
    .B1(_00775_),
    .Y(_00777_));
 sky130_fd_sc_hd__xor2_1 _07364_ (.A(_00771_),
    .B(_00777_),
    .X(net81));
 sky130_fd_sc_hd__nor2_1 _07365_ (.A(_00659_),
    .B(_00661_),
    .Y(_00779_));
 sky130_fd_sc_hd__a31o_1 _07366_ (.A1(net12),
    .A2(net48),
    .A3(_00649_),
    .B1(_00646_),
    .X(_00780_));
 sky130_fd_sc_hd__a22o_1 _07367_ (.A1(net12),
    .A2(net49),
    .B1(net50),
    .B2(net1),
    .X(_00781_));
 sky130_fd_sc_hd__and4_1 _07368_ (.A(net12),
    .B(net1),
    .C(net49),
    .D(net50),
    .X(_00782_));
 sky130_fd_sc_hd__inv_2 _07369_ (.A(_00782_),
    .Y(_00783_));
 sky130_fd_sc_hd__and3_1 _07370_ (.A(_00780_),
    .B(_00781_),
    .C(_00783_),
    .X(_00784_));
 sky130_fd_sc_hd__a21oi_1 _07371_ (.A1(_00781_),
    .A2(_00783_),
    .B1(_00780_),
    .Y(_00785_));
 sky130_fd_sc_hd__nor2_1 _07372_ (.A(_00784_),
    .B(_00785_),
    .Y(_00786_));
 sky130_fd_sc_hd__or3_1 _07373_ (.A(_00779_),
    .B(_00784_),
    .C(_00785_),
    .X(_00787_));
 sky130_fd_sc_hd__xnor2_1 _07374_ (.A(_00779_),
    .B(_00786_),
    .Y(_00788_));
 sky130_fd_sc_hd__nand2_1 _07375_ (.A(_00635_),
    .B(_00788_),
    .Y(_00790_));
 sky130_fd_sc_hd__xnor2_1 _07376_ (.A(_00635_),
    .B(_00788_),
    .Y(_00791_));
 sky130_fd_sc_hd__nor2_1 _07377_ (.A(_00639_),
    .B(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hd__xor2_1 _07378_ (.A(_00639_),
    .B(_00791_),
    .X(_00793_));
 sky130_fd_sc_hd__nor3_1 _07379_ (.A(_00684_),
    .B(_00686_),
    .C(_00793_),
    .Y(_00794_));
 sky130_fd_sc_hd__o21a_1 _07380_ (.A1(_00684_),
    .A2(_00686_),
    .B1(_00793_),
    .X(_00795_));
 sky130_fd_sc_hd__nor2_1 _07381_ (.A(_00794_),
    .B(_00795_),
    .Y(_00796_));
 sky130_fd_sc_hd__and2_1 _07382_ (.A(_00642_),
    .B(_00796_),
    .X(_00797_));
 sky130_fd_sc_hd__xnor2_1 _07383_ (.A(_00642_),
    .B(_00796_),
    .Y(_00798_));
 sky130_fd_sc_hd__nand2_1 _07384_ (.A(net23),
    .B(net48),
    .Y(_00799_));
 sky130_fd_sc_hd__and4_1 _07385_ (.A(net27),
    .B(net26),
    .C(net46),
    .D(net47),
    .X(_00801_));
 sky130_fd_sc_hd__a22o_1 _07386_ (.A1(net27),
    .A2(net46),
    .B1(net47),
    .B2(net26),
    .X(_00802_));
 sky130_fd_sc_hd__and2b_1 _07387_ (.A_N(_00801_),
    .B(_00802_),
    .X(_00803_));
 sky130_fd_sc_hd__xnor2_1 _07388_ (.A(_00799_),
    .B(_00803_),
    .Y(_00804_));
 sky130_fd_sc_hd__nand2_1 _07389_ (.A(net28),
    .B(net45),
    .Y(_00805_));
 sky130_fd_sc_hd__and4_1 _07390_ (.A(net29),
    .B(net30),
    .C(net42),
    .D(net43),
    .X(_00806_));
 sky130_fd_sc_hd__a22oi_2 _07391_ (.A1(net30),
    .A2(net42),
    .B1(net43),
    .B2(net29),
    .Y(_00807_));
 sky130_fd_sc_hd__or3_1 _07392_ (.A(_00805_),
    .B(_00806_),
    .C(_00807_),
    .X(_00808_));
 sky130_fd_sc_hd__o21ai_1 _07393_ (.A1(_00806_),
    .A2(_00807_),
    .B1(_00805_),
    .Y(_00809_));
 sky130_fd_sc_hd__o21bai_1 _07394_ (.A1(_00653_),
    .A2(_00654_),
    .B1_N(_00652_),
    .Y(_00810_));
 sky130_fd_sc_hd__and3_1 _07395_ (.A(_00808_),
    .B(_00809_),
    .C(_00810_),
    .X(_00812_));
 sky130_fd_sc_hd__a21o_1 _07396_ (.A1(_00808_),
    .A2(_00809_),
    .B1(_00810_),
    .X(_00813_));
 sky130_fd_sc_hd__and2b_1 _07397_ (.A_N(_00812_),
    .B(_00813_),
    .X(_00814_));
 sky130_fd_sc_hd__xnor2_1 _07398_ (.A(_00804_),
    .B(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_1 _07399_ (.A(_00666_),
    .B(_00670_),
    .Y(_00816_));
 sky130_fd_sc_hd__a31o_1 _07400_ (.A1(net2),
    .A2(net38),
    .A3(_00690_),
    .B1(_00689_),
    .X(_00817_));
 sky130_fd_sc_hd__nand4_2 _07401_ (.A(net2),
    .B(net32),
    .C(net39),
    .D(net40),
    .Y(_00818_));
 sky130_fd_sc_hd__a22o_1 _07402_ (.A1(net2),
    .A2(net39),
    .B1(net40),
    .B2(net32),
    .X(_00819_));
 sky130_fd_sc_hd__nand4_2 _07403_ (.A(net31),
    .B(net41),
    .C(_00818_),
    .D(_00819_),
    .Y(_00820_));
 sky130_fd_sc_hd__a22o_1 _07404_ (.A1(net31),
    .A2(net41),
    .B1(_00818_),
    .B2(_00819_),
    .X(_00821_));
 sky130_fd_sc_hd__nand3_2 _07405_ (.A(_00817_),
    .B(_00820_),
    .C(_00821_),
    .Y(_00823_));
 sky130_fd_sc_hd__a21o_1 _07406_ (.A1(_00820_),
    .A2(_00821_),
    .B1(_00817_),
    .X(_00824_));
 sky130_fd_sc_hd__nand3_2 _07407_ (.A(_00816_),
    .B(_00823_),
    .C(_00824_),
    .Y(_00825_));
 sky130_fd_sc_hd__a21o_1 _07408_ (.A1(_00823_),
    .A2(_00824_),
    .B1(_00816_),
    .X(_00826_));
 sky130_fd_sc_hd__a21bo_1 _07409_ (.A1(_00664_),
    .A2(_00673_),
    .B1_N(_00672_),
    .X(_00827_));
 sky130_fd_sc_hd__and3_1 _07410_ (.A(_00825_),
    .B(_00826_),
    .C(_00827_),
    .X(_00828_));
 sky130_fd_sc_hd__nand3_1 _07411_ (.A(_00825_),
    .B(_00826_),
    .C(_00827_),
    .Y(_00829_));
 sky130_fd_sc_hd__a21oi_1 _07412_ (.A1(_00825_),
    .A2(_00826_),
    .B1(_00827_),
    .Y(_00830_));
 sky130_fd_sc_hd__or3_2 _07413_ (.A(_00815_),
    .B(_00828_),
    .C(_00830_),
    .X(_00831_));
 sky130_fd_sc_hd__o21ai_1 _07414_ (.A1(_00828_),
    .A2(_00830_),
    .B1(_00815_),
    .Y(_00832_));
 sky130_fd_sc_hd__o211a_1 _07415_ (.A1(_00706_),
    .A2(_00708_),
    .B1(_00831_),
    .C1(_00832_),
    .X(_00834_));
 sky130_fd_sc_hd__a211oi_1 _07416_ (.A1(_00831_),
    .A2(_00832_),
    .B1(_00706_),
    .C1(_00708_),
    .Y(_00835_));
 sky130_fd_sc_hd__a211oi_1 _07417_ (.A1(_00678_),
    .A2(_00682_),
    .B1(_00834_),
    .C1(_00835_),
    .Y(_00836_));
 sky130_fd_sc_hd__o211a_1 _07418_ (.A1(_00834_),
    .A2(_00835_),
    .B1(_00678_),
    .C1(_00682_),
    .X(_00837_));
 sky130_fd_sc_hd__nand2_1 _07419_ (.A(net3),
    .B(net38),
    .Y(_00838_));
 sky130_fd_sc_hd__and4_1 _07420_ (.A(net4),
    .B(net36),
    .C(net5),
    .D(net37),
    .X(_00839_));
 sky130_fd_sc_hd__a22oi_1 _07421_ (.A1(net36),
    .A2(net5),
    .B1(net37),
    .B2(net4),
    .Y(_00840_));
 sky130_fd_sc_hd__nor2_1 _07422_ (.A(_00839_),
    .B(_00840_),
    .Y(_00841_));
 sky130_fd_sc_hd__xnor2_1 _07423_ (.A(_00838_),
    .B(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__and4_1 _07424_ (.A(net64),
    .B(net34),
    .C(net7),
    .D(net8),
    .X(_00843_));
 sky130_fd_sc_hd__a22oi_1 _07425_ (.A1(net34),
    .A2(net7),
    .B1(net8),
    .B2(net64),
    .Y(_00845_));
 sky130_fd_sc_hd__and4bb_1 _07426_ (.A_N(_00843_),
    .B_N(_00845_),
    .C(net35),
    .D(net6),
    .X(_00846_));
 sky130_fd_sc_hd__o2bb2a_1 _07427_ (.A1_N(net35),
    .A2_N(net6),
    .B1(_00843_),
    .B2(_00845_),
    .X(_00847_));
 sky130_fd_sc_hd__nor2_1 _07428_ (.A(_00846_),
    .B(_00847_),
    .Y(_00848_));
 sky130_fd_sc_hd__nand2_1 _07429_ (.A(_00695_),
    .B(_00698_),
    .Y(_00849_));
 sky130_fd_sc_hd__and2_1 _07430_ (.A(_00848_),
    .B(_00849_),
    .X(_00850_));
 sky130_fd_sc_hd__xor2_1 _07431_ (.A(_00848_),
    .B(_00849_),
    .X(_00851_));
 sky130_fd_sc_hd__and2_1 _07432_ (.A(_00842_),
    .B(_00851_),
    .X(_00852_));
 sky130_fd_sc_hd__xnor2_1 _07433_ (.A(_00842_),
    .B(_00851_),
    .Y(_00853_));
 sky130_fd_sc_hd__a21oi_2 _07434_ (.A1(_00718_),
    .A2(_00720_),
    .B1(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__inv_2 _07435_ (.A(_00854_),
    .Y(_00855_));
 sky130_fd_sc_hd__and3_1 _07436_ (.A(_00718_),
    .B(_00720_),
    .C(_00853_),
    .X(_00856_));
 sky130_fd_sc_hd__a211oi_1 _07437_ (.A1(_00701_),
    .A2(_00704_),
    .B1(_00854_),
    .C1(_00856_),
    .Y(_00857_));
 sky130_fd_sc_hd__a211o_1 _07438_ (.A1(_00701_),
    .A2(_00704_),
    .B1(_00854_),
    .C1(_00856_),
    .X(_00858_));
 sky130_fd_sc_hd__o211a_1 _07439_ (.A1(_00854_),
    .A2(_00856_),
    .B1(_00701_),
    .C1(_00704_),
    .X(_00859_));
 sky130_fd_sc_hd__o21ba_1 _07440_ (.A1(_00714_),
    .A2(_00716_),
    .B1_N(_00712_),
    .X(_00860_));
 sky130_fd_sc_hd__o21ba_1 _07441_ (.A1(_00723_),
    .A2(_00726_),
    .B1_N(_00722_),
    .X(_00861_));
 sky130_fd_sc_hd__nand2_1 _07442_ (.A(net63),
    .B(net9),
    .Y(_00862_));
 sky130_fd_sc_hd__and4_1 _07443_ (.A(net61),
    .B(net62),
    .C(net10),
    .D(net11),
    .X(_00863_));
 sky130_fd_sc_hd__a22oi_1 _07444_ (.A1(net62),
    .A2(net10),
    .B1(net11),
    .B2(net61),
    .Y(_00864_));
 sky130_fd_sc_hd__nor2_1 _07445_ (.A(_00863_),
    .B(_00864_),
    .Y(_00866_));
 sky130_fd_sc_hd__xnor2_1 _07446_ (.A(_00862_),
    .B(_00866_),
    .Y(_00867_));
 sky130_fd_sc_hd__nand2b_1 _07447_ (.A_N(_00861_),
    .B(_00867_),
    .Y(_00868_));
 sky130_fd_sc_hd__xnor2_1 _07448_ (.A(_00861_),
    .B(_00867_),
    .Y(_00869_));
 sky130_fd_sc_hd__nand2b_1 _07449_ (.A_N(_00860_),
    .B(_00869_),
    .Y(_00870_));
 sky130_fd_sc_hd__xnor2_1 _07450_ (.A(_00860_),
    .B(_00869_),
    .Y(_00871_));
 sky130_fd_sc_hd__nand2_1 _07451_ (.A(net60),
    .B(net13),
    .Y(_00872_));
 sky130_fd_sc_hd__and4_1 _07452_ (.A(net58),
    .B(net59),
    .C(net14),
    .D(net15),
    .X(_00873_));
 sky130_fd_sc_hd__a22oi_1 _07453_ (.A1(net59),
    .A2(net14),
    .B1(net15),
    .B2(net58),
    .Y(_00874_));
 sky130_fd_sc_hd__nor2_1 _07454_ (.A(_00873_),
    .B(_00874_),
    .Y(_00875_));
 sky130_fd_sc_hd__xnor2_1 _07455_ (.A(_00872_),
    .B(_00875_),
    .Y(_00877_));
 sky130_fd_sc_hd__and2_1 _07456_ (.A(net55),
    .B(net16),
    .X(_00878_));
 sky130_fd_sc_hd__nand4_1 _07457_ (.A(net33),
    .B(net44),
    .C(net17),
    .D(net18),
    .Y(_00879_));
 sky130_fd_sc_hd__a22o_1 _07458_ (.A1(net44),
    .A2(net17),
    .B1(net18),
    .B2(net33),
    .X(_00880_));
 sky130_fd_sc_hd__nand3_1 _07459_ (.A(_00878_),
    .B(_00879_),
    .C(_00880_),
    .Y(_00881_));
 sky130_fd_sc_hd__a21o_1 _07460_ (.A1(_00879_),
    .A2(_00880_),
    .B1(_00878_),
    .X(_00882_));
 sky130_fd_sc_hd__o21bai_1 _07461_ (.A1(_00728_),
    .A2(_00730_),
    .B1_N(_00729_),
    .Y(_00883_));
 sky130_fd_sc_hd__nand3_1 _07462_ (.A(_00881_),
    .B(_00882_),
    .C(_00883_),
    .Y(_00884_));
 sky130_fd_sc_hd__a21o_1 _07463_ (.A1(_00881_),
    .A2(_00882_),
    .B1(_00883_),
    .X(_00885_));
 sky130_fd_sc_hd__nand3_1 _07464_ (.A(_00877_),
    .B(_00884_),
    .C(_00885_),
    .Y(_00886_));
 sky130_fd_sc_hd__a21o_1 _07465_ (.A1(_00884_),
    .A2(_00885_),
    .B1(_00877_),
    .X(_00888_));
 sky130_fd_sc_hd__a21bo_1 _07466_ (.A1(_00727_),
    .A2(_00736_),
    .B1_N(_00734_),
    .X(_00889_));
 sky130_fd_sc_hd__nand3_2 _07467_ (.A(_00886_),
    .B(_00888_),
    .C(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__a21o_1 _07468_ (.A1(_00886_),
    .A2(_00888_),
    .B1(_00889_),
    .X(_00891_));
 sky130_fd_sc_hd__and3_1 _07469_ (.A(_00871_),
    .B(_00890_),
    .C(_00891_),
    .X(_00892_));
 sky130_fd_sc_hd__nand3_1 _07470_ (.A(_00871_),
    .B(_00890_),
    .C(_00891_),
    .Y(_00893_));
 sky130_fd_sc_hd__a21oi_2 _07471_ (.A1(_00890_),
    .A2(_00891_),
    .B1(_00871_),
    .Y(_00894_));
 sky130_fd_sc_hd__a211oi_4 _07472_ (.A1(_00740_),
    .A2(_00743_),
    .B1(_00892_),
    .C1(_00894_),
    .Y(_00895_));
 sky130_fd_sc_hd__o211a_1 _07473_ (.A1(_00892_),
    .A2(_00894_),
    .B1(_00740_),
    .C1(_00743_),
    .X(_00896_));
 sky130_fd_sc_hd__nor4_2 _07474_ (.A(_00857_),
    .B(_00859_),
    .C(_00895_),
    .D(_00896_),
    .Y(_00897_));
 sky130_fd_sc_hd__o22a_1 _07475_ (.A1(_00857_),
    .A2(_00859_),
    .B1(_00895_),
    .B2(_00896_),
    .X(_00899_));
 sky130_fd_sc_hd__a211o_1 _07476_ (.A1(_00745_),
    .A2(_00748_),
    .B1(_00897_),
    .C1(_00899_),
    .X(_00900_));
 sky130_fd_sc_hd__o211ai_1 _07477_ (.A1(_00897_),
    .A2(_00899_),
    .B1(_00745_),
    .C1(_00748_),
    .Y(_00901_));
 sky130_fd_sc_hd__or4bb_2 _07478_ (.A(_00836_),
    .B(_00837_),
    .C_N(_00900_),
    .D_N(_00901_),
    .X(_00902_));
 sky130_fd_sc_hd__a2bb2o_1 _07479_ (.A1_N(_00836_),
    .A2_N(_00837_),
    .B1(_00900_),
    .B2(_00901_),
    .X(_00903_));
 sky130_fd_sc_hd__o211a_2 _07480_ (.A1(_00750_),
    .A2(_00752_),
    .B1(_00902_),
    .C1(_00903_),
    .X(_00904_));
 sky130_fd_sc_hd__a211oi_1 _07481_ (.A1(_00902_),
    .A2(_00903_),
    .B1(_00750_),
    .C1(_00752_),
    .Y(_00905_));
 sky130_fd_sc_hd__nor3_1 _07482_ (.A(_00798_),
    .B(_00904_),
    .C(_00905_),
    .Y(_00906_));
 sky130_fd_sc_hd__or3_1 _07483_ (.A(_00798_),
    .B(_00904_),
    .C(_00905_),
    .X(_00907_));
 sky130_fd_sc_hd__o21ai_1 _07484_ (.A1(_00904_),
    .A2(_00905_),
    .B1(_00798_),
    .Y(_00908_));
 sky130_fd_sc_hd__o211a_1 _07485_ (.A1(_00754_),
    .A2(_00756_),
    .B1(_00907_),
    .C1(_00908_),
    .X(_00910_));
 sky130_fd_sc_hd__o211ai_1 _07486_ (.A1(_00754_),
    .A2(_00756_),
    .B1(_00907_),
    .C1(_00908_),
    .Y(_00911_));
 sky130_fd_sc_hd__a211oi_1 _07487_ (.A1(_00907_),
    .A2(_00908_),
    .B1(_00754_),
    .C1(_00756_),
    .Y(_00912_));
 sky130_fd_sc_hd__or3_2 _07488_ (.A(_00644_),
    .B(_00910_),
    .C(_00912_),
    .X(_00913_));
 sky130_fd_sc_hd__o21ai_1 _07489_ (.A1(_00910_),
    .A2(_00912_),
    .B1(_00644_),
    .Y(_00914_));
 sky130_fd_sc_hd__o211ai_2 _07490_ (.A1(_00760_),
    .A2(_00763_),
    .B1(_00913_),
    .C1(_00914_),
    .Y(_00915_));
 sky130_fd_sc_hd__a211o_1 _07491_ (.A1(_00913_),
    .A2(_00914_),
    .B1(_00760_),
    .C1(_00763_),
    .X(_00916_));
 sky130_fd_sc_hd__a21oi_1 _07492_ (.A1(_00915_),
    .A2(_00916_),
    .B1(_00766_),
    .Y(_00917_));
 sky130_fd_sc_hd__and3_1 _07493_ (.A(_00766_),
    .B(_00915_),
    .C(_00916_),
    .X(_00918_));
 sky130_fd_sc_hd__nor2_1 _07494_ (.A(_00917_),
    .B(_00918_),
    .Y(_00919_));
 sky130_fd_sc_hd__o21ba_1 _07495_ (.A1(_00771_),
    .A2(_00777_),
    .B1_N(_00770_),
    .X(_00921_));
 sky130_fd_sc_hd__xnor2_1 _07496_ (.A(_00919_),
    .B(_00921_),
    .Y(net82));
 sky130_fd_sc_hd__or2_1 _07497_ (.A(_00834_),
    .B(_00836_),
    .X(_00922_));
 sky130_fd_sc_hd__a21oi_1 _07498_ (.A1(_00804_),
    .A2(_00813_),
    .B1(_00812_),
    .Y(_00923_));
 sky130_fd_sc_hd__a31o_1 _07499_ (.A1(net23),
    .A2(net48),
    .A3(_00802_),
    .B1(_00801_),
    .X(_00924_));
 sky130_fd_sc_hd__nand4_1 _07500_ (.A(net23),
    .B(net12),
    .C(net49),
    .D(net50),
    .Y(_00925_));
 sky130_fd_sc_hd__a22o_1 _07501_ (.A1(net23),
    .A2(net49),
    .B1(net50),
    .B2(net12),
    .X(_00926_));
 sky130_fd_sc_hd__nand2_1 _07502_ (.A(net1),
    .B(net51),
    .Y(_00927_));
 sky130_fd_sc_hd__nand3b_1 _07503_ (.A_N(_00927_),
    .B(_00926_),
    .C(_00925_),
    .Y(_00928_));
 sky130_fd_sc_hd__a21bo_1 _07504_ (.A1(_00925_),
    .A2(_00926_),
    .B1_N(_00927_),
    .X(_00929_));
 sky130_fd_sc_hd__and3_1 _07505_ (.A(_00924_),
    .B(_00928_),
    .C(_00929_),
    .X(_00931_));
 sky130_fd_sc_hd__a21o_1 _07506_ (.A1(_00928_),
    .A2(_00929_),
    .B1(_00924_),
    .X(_00932_));
 sky130_fd_sc_hd__and2b_1 _07507_ (.A_N(_00931_),
    .B(_00932_),
    .X(_00933_));
 sky130_fd_sc_hd__xnor2_1 _07508_ (.A(_00782_),
    .B(_00933_),
    .Y(_00934_));
 sky130_fd_sc_hd__nor2_1 _07509_ (.A(_00923_),
    .B(_00934_),
    .Y(_00935_));
 sky130_fd_sc_hd__xor2_1 _07510_ (.A(_00923_),
    .B(_00934_),
    .X(_00936_));
 sky130_fd_sc_hd__xnor2_1 _07511_ (.A(_00784_),
    .B(_00936_),
    .Y(_00937_));
 sky130_fd_sc_hd__a21o_1 _07512_ (.A1(_00787_),
    .A2(_00790_),
    .B1(_00937_),
    .X(_00938_));
 sky130_fd_sc_hd__nand3_1 _07513_ (.A(_00787_),
    .B(_00790_),
    .C(_00937_),
    .Y(_00939_));
 sky130_fd_sc_hd__nand2_1 _07514_ (.A(_00938_),
    .B(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand2b_1 _07515_ (.A_N(_00940_),
    .B(_00922_),
    .Y(_00942_));
 sky130_fd_sc_hd__xnor2_1 _07516_ (.A(_00922_),
    .B(_00940_),
    .Y(_00943_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(_00792_),
    .B(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__xnor2_1 _07518_ (.A(_00792_),
    .B(_00943_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand2_1 _07519_ (.A(net26),
    .B(net48),
    .Y(_00946_));
 sky130_fd_sc_hd__and4_1 _07520_ (.A(net28),
    .B(net27),
    .C(net46),
    .D(net47),
    .X(_00947_));
 sky130_fd_sc_hd__a22oi_1 _07521_ (.A1(net28),
    .A2(net46),
    .B1(net47),
    .B2(net27),
    .Y(_00948_));
 sky130_fd_sc_hd__nor2_1 _07522_ (.A(_00947_),
    .B(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__xnor2_1 _07523_ (.A(_00946_),
    .B(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__and4_1 _07524_ (.A(net30),
    .B(net31),
    .C(net42),
    .D(net43),
    .X(_00951_));
 sky130_fd_sc_hd__a22oi_1 _07525_ (.A1(net31),
    .A2(net42),
    .B1(net43),
    .B2(net30),
    .Y(_00953_));
 sky130_fd_sc_hd__and4bb_1 _07526_ (.A_N(_00951_),
    .B_N(_00953_),
    .C(net29),
    .D(net45),
    .X(_00954_));
 sky130_fd_sc_hd__o2bb2a_1 _07527_ (.A1_N(net29),
    .A2_N(net45),
    .B1(_00951_),
    .B2(_00953_),
    .X(_00955_));
 sky130_fd_sc_hd__o21ba_1 _07528_ (.A1(_00805_),
    .A2(_00807_),
    .B1_N(_00806_),
    .X(_00956_));
 sky130_fd_sc_hd__nor3_1 _07529_ (.A(_00954_),
    .B(_00955_),
    .C(_00956_),
    .Y(_00957_));
 sky130_fd_sc_hd__o21a_1 _07530_ (.A1(_00954_),
    .A2(_00955_),
    .B1(_00956_),
    .X(_00958_));
 sky130_fd_sc_hd__nor2_1 _07531_ (.A(_00957_),
    .B(_00958_),
    .Y(_00959_));
 sky130_fd_sc_hd__xnor2_1 _07532_ (.A(_00950_),
    .B(_00959_),
    .Y(_00960_));
 sky130_fd_sc_hd__nand2_1 _07533_ (.A(_00818_),
    .B(_00820_),
    .Y(_00961_));
 sky130_fd_sc_hd__o21ba_1 _07534_ (.A1(_00838_),
    .A2(_00840_),
    .B1_N(_00839_),
    .X(_00962_));
 sky130_fd_sc_hd__nand2_1 _07535_ (.A(net32),
    .B(net41),
    .Y(_00963_));
 sky130_fd_sc_hd__and4_1 _07536_ (.A(net2),
    .B(net3),
    .C(net39),
    .D(net40),
    .X(_00964_));
 sky130_fd_sc_hd__a22oi_1 _07537_ (.A1(net3),
    .A2(net39),
    .B1(net40),
    .B2(net2),
    .Y(_00965_));
 sky130_fd_sc_hd__nor2_1 _07538_ (.A(_00964_),
    .B(_00965_),
    .Y(_00966_));
 sky130_fd_sc_hd__xnor2_1 _07539_ (.A(_00963_),
    .B(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__nand2b_1 _07540_ (.A_N(_00962_),
    .B(_00967_),
    .Y(_00968_));
 sky130_fd_sc_hd__xnor2_1 _07541_ (.A(_00962_),
    .B(_00967_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_1 _07542_ (.A(_00961_),
    .B(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__xnor2_1 _07543_ (.A(_00961_),
    .B(_00969_),
    .Y(_00971_));
 sky130_fd_sc_hd__a21oi_2 _07544_ (.A1(_00823_),
    .A2(_00825_),
    .B1(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__inv_2 _07545_ (.A(_00972_),
    .Y(_00974_));
 sky130_fd_sc_hd__and3_1 _07546_ (.A(_00823_),
    .B(_00825_),
    .C(_00971_),
    .X(_00975_));
 sky130_fd_sc_hd__nor3_2 _07547_ (.A(_00960_),
    .B(_00972_),
    .C(_00975_),
    .Y(_00976_));
 sky130_fd_sc_hd__inv_2 _07548_ (.A(_00976_),
    .Y(_00977_));
 sky130_fd_sc_hd__o21a_1 _07549_ (.A1(_00972_),
    .A2(_00975_),
    .B1(_00960_),
    .X(_00978_));
 sky130_fd_sc_hd__a211oi_4 _07550_ (.A1(_00855_),
    .A2(_00858_),
    .B1(_00976_),
    .C1(_00978_),
    .Y(_00979_));
 sky130_fd_sc_hd__o211a_1 _07551_ (.A1(_00976_),
    .A2(_00978_),
    .B1(_00855_),
    .C1(_00858_),
    .X(_00980_));
 sky130_fd_sc_hd__a211oi_4 _07552_ (.A1(_00829_),
    .A2(_00831_),
    .B1(_00979_),
    .C1(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__o211a_1 _07553_ (.A1(_00979_),
    .A2(_00980_),
    .B1(_00829_),
    .C1(_00831_),
    .X(_00982_));
 sky130_fd_sc_hd__nand2_1 _07554_ (.A(net4),
    .B(net38),
    .Y(_00983_));
 sky130_fd_sc_hd__and4_1 _07555_ (.A(net36),
    .B(net5),
    .C(net37),
    .D(net6),
    .X(_00985_));
 sky130_fd_sc_hd__a22oi_1 _07556_ (.A1(net5),
    .A2(net37),
    .B1(net6),
    .B2(net36),
    .Y(_00986_));
 sky130_fd_sc_hd__nor2_1 _07557_ (.A(_00985_),
    .B(_00986_),
    .Y(_00987_));
 sky130_fd_sc_hd__xnor2_1 _07558_ (.A(_00983_),
    .B(_00987_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _07559_ (.A(net35),
    .B(net7),
    .Y(_00989_));
 sky130_fd_sc_hd__and4_1 _07560_ (.A(net64),
    .B(net34),
    .C(net8),
    .D(net9),
    .X(_00990_));
 sky130_fd_sc_hd__a22oi_1 _07561_ (.A1(net34),
    .A2(net8),
    .B1(net9),
    .B2(net64),
    .Y(_00991_));
 sky130_fd_sc_hd__nor2_1 _07562_ (.A(_00990_),
    .B(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__xnor2_1 _07563_ (.A(_00989_),
    .B(_00992_),
    .Y(_00993_));
 sky130_fd_sc_hd__nor2_1 _07564_ (.A(_00843_),
    .B(_00846_),
    .Y(_00994_));
 sky130_fd_sc_hd__and2b_1 _07565_ (.A_N(_00994_),
    .B(_00993_),
    .X(_00996_));
 sky130_fd_sc_hd__xnor2_1 _07566_ (.A(_00993_),
    .B(_00994_),
    .Y(_00997_));
 sky130_fd_sc_hd__and2_1 _07567_ (.A(_00988_),
    .B(_00997_),
    .X(_00998_));
 sky130_fd_sc_hd__xnor2_1 _07568_ (.A(_00988_),
    .B(_00997_),
    .Y(_00999_));
 sky130_fd_sc_hd__a21oi_1 _07569_ (.A1(_00868_),
    .A2(_00870_),
    .B1(_00999_),
    .Y(_01000_));
 sky130_fd_sc_hd__a21o_1 _07570_ (.A1(_00868_),
    .A2(_00870_),
    .B1(_00999_),
    .X(_01001_));
 sky130_fd_sc_hd__nand3_1 _07571_ (.A(_00868_),
    .B(_00870_),
    .C(_00999_),
    .Y(_01002_));
 sky130_fd_sc_hd__o211a_1 _07572_ (.A1(_00850_),
    .A2(_00852_),
    .B1(_01001_),
    .C1(_01002_),
    .X(_01003_));
 sky130_fd_sc_hd__a211oi_1 _07573_ (.A1(_01001_),
    .A2(_01002_),
    .B1(_00850_),
    .C1(_00852_),
    .Y(_01004_));
 sky130_fd_sc_hd__o21ba_1 _07574_ (.A1(_00862_),
    .A2(_00864_),
    .B1_N(_00863_),
    .X(_01005_));
 sky130_fd_sc_hd__o21ba_1 _07575_ (.A1(_00872_),
    .A2(_00874_),
    .B1_N(_00873_),
    .X(_01007_));
 sky130_fd_sc_hd__nand2_1 _07576_ (.A(net63),
    .B(net10),
    .Y(_01008_));
 sky130_fd_sc_hd__and4_1 _07577_ (.A(net61),
    .B(net62),
    .C(net11),
    .D(net13),
    .X(_01009_));
 sky130_fd_sc_hd__a22oi_1 _07578_ (.A1(net62),
    .A2(net11),
    .B1(net13),
    .B2(net61),
    .Y(_01010_));
 sky130_fd_sc_hd__nor2_1 _07579_ (.A(_01009_),
    .B(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__xnor2_1 _07580_ (.A(_01008_),
    .B(_01011_),
    .Y(_01012_));
 sky130_fd_sc_hd__nand2b_1 _07581_ (.A_N(_01007_),
    .B(_01012_),
    .Y(_01013_));
 sky130_fd_sc_hd__xnor2_1 _07582_ (.A(_01007_),
    .B(_01012_),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2b_1 _07583_ (.A_N(_01005_),
    .B(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hd__xnor2_1 _07584_ (.A(_01005_),
    .B(_01014_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_1 _07585_ (.A(net60),
    .B(net14),
    .Y(_01018_));
 sky130_fd_sc_hd__and4_1 _07586_ (.A(net58),
    .B(net59),
    .C(net15),
    .D(net16),
    .X(_01019_));
 sky130_fd_sc_hd__a22oi_1 _07587_ (.A1(net59),
    .A2(net15),
    .B1(net16),
    .B2(net58),
    .Y(_01020_));
 sky130_fd_sc_hd__nor2_1 _07588_ (.A(_01019_),
    .B(_01020_),
    .Y(_01021_));
 sky130_fd_sc_hd__xnor2_1 _07589_ (.A(_01018_),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__nand2_1 _07590_ (.A(net55),
    .B(net17),
    .Y(_01023_));
 sky130_fd_sc_hd__and4_1 _07591_ (.A(net33),
    .B(net44),
    .C(net18),
    .D(net19),
    .X(_01024_));
 sky130_fd_sc_hd__a22oi_2 _07592_ (.A1(net44),
    .A2(net18),
    .B1(net19),
    .B2(net33),
    .Y(_01025_));
 sky130_fd_sc_hd__or3_1 _07593_ (.A(_01023_),
    .B(_01024_),
    .C(_01025_),
    .X(_01026_));
 sky130_fd_sc_hd__o21ai_1 _07594_ (.A1(_01024_),
    .A2(_01025_),
    .B1(_01023_),
    .Y(_01027_));
 sky130_fd_sc_hd__a21bo_1 _07595_ (.A1(_00878_),
    .A2(_00880_),
    .B1_N(_00879_),
    .X(_01029_));
 sky130_fd_sc_hd__nand3_1 _07596_ (.A(_01026_),
    .B(_01027_),
    .C(_01029_),
    .Y(_01030_));
 sky130_fd_sc_hd__a21o_1 _07597_ (.A1(_01026_),
    .A2(_01027_),
    .B1(_01029_),
    .X(_01031_));
 sky130_fd_sc_hd__nand3_1 _07598_ (.A(_01022_),
    .B(_01030_),
    .C(_01031_),
    .Y(_01032_));
 sky130_fd_sc_hd__a21o_1 _07599_ (.A1(_01030_),
    .A2(_01031_),
    .B1(_01022_),
    .X(_01033_));
 sky130_fd_sc_hd__a21bo_1 _07600_ (.A1(_00877_),
    .A2(_00885_),
    .B1_N(_00884_),
    .X(_01034_));
 sky130_fd_sc_hd__nand3_4 _07601_ (.A(_01032_),
    .B(_01033_),
    .C(_01034_),
    .Y(_01035_));
 sky130_fd_sc_hd__a21o_1 _07602_ (.A1(_01032_),
    .A2(_01033_),
    .B1(_01034_),
    .X(_01036_));
 sky130_fd_sc_hd__and3_1 _07603_ (.A(_01016_),
    .B(_01035_),
    .C(_01036_),
    .X(_01037_));
 sky130_fd_sc_hd__nand3_2 _07604_ (.A(_01016_),
    .B(_01035_),
    .C(_01036_),
    .Y(_01038_));
 sky130_fd_sc_hd__a21oi_1 _07605_ (.A1(_01035_),
    .A2(_01036_),
    .B1(_01016_),
    .Y(_01040_));
 sky130_fd_sc_hd__a211o_1 _07606_ (.A1(_00890_),
    .A2(_00893_),
    .B1(_01037_),
    .C1(_01040_),
    .X(_01041_));
 sky130_fd_sc_hd__o211ai_1 _07607_ (.A1(_01037_),
    .A2(_01040_),
    .B1(_00890_),
    .C1(_00893_),
    .Y(_01042_));
 sky130_fd_sc_hd__or4bb_2 _07608_ (.A(_01003_),
    .B(_01004_),
    .C_N(_01041_),
    .D_N(_01042_),
    .X(_01043_));
 sky130_fd_sc_hd__a2bb2o_1 _07609_ (.A1_N(_01003_),
    .A2_N(_01004_),
    .B1(_01041_),
    .B2(_01042_),
    .X(_01044_));
 sky130_fd_sc_hd__o211a_2 _07610_ (.A1(_00895_),
    .A2(_00897_),
    .B1(_01043_),
    .C1(_01044_),
    .X(_01045_));
 sky130_fd_sc_hd__a211oi_2 _07611_ (.A1(_01043_),
    .A2(_01044_),
    .B1(_00895_),
    .C1(_00897_),
    .Y(_01046_));
 sky130_fd_sc_hd__nor4_4 _07612_ (.A(_00981_),
    .B(_00982_),
    .C(_01045_),
    .D(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__o22a_1 _07613_ (.A1(_00981_),
    .A2(_00982_),
    .B1(_01045_),
    .B2(_01046_),
    .X(_01048_));
 sky130_fd_sc_hd__a211oi_4 _07614_ (.A1(_00900_),
    .A2(_00902_),
    .B1(_01047_),
    .C1(_01048_),
    .Y(_01049_));
 sky130_fd_sc_hd__o211a_1 _07615_ (.A1(_01047_),
    .A2(_01048_),
    .B1(_00900_),
    .C1(_00902_),
    .X(_01051_));
 sky130_fd_sc_hd__nor3_1 _07616_ (.A(_00945_),
    .B(_01049_),
    .C(_01051_),
    .Y(_01052_));
 sky130_fd_sc_hd__or3_2 _07617_ (.A(_00945_),
    .B(_01049_),
    .C(_01051_),
    .X(_01053_));
 sky130_fd_sc_hd__o21ai_2 _07618_ (.A1(_01049_),
    .A2(_01051_),
    .B1(_00945_),
    .Y(_01054_));
 sky130_fd_sc_hd__o211ai_4 _07619_ (.A1(_00904_),
    .A2(_00906_),
    .B1(_01053_),
    .C1(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hd__a211o_1 _07620_ (.A1(_01053_),
    .A2(_01054_),
    .B1(_00904_),
    .C1(_00906_),
    .X(_01056_));
 sky130_fd_sc_hd__o211a_1 _07621_ (.A1(_00795_),
    .A2(_00797_),
    .B1(_01055_),
    .C1(_01056_),
    .X(_01057_));
 sky130_fd_sc_hd__o211ai_2 _07622_ (.A1(_00795_),
    .A2(_00797_),
    .B1(_01055_),
    .C1(_01056_),
    .Y(_01058_));
 sky130_fd_sc_hd__a211oi_1 _07623_ (.A1(_01055_),
    .A2(_01056_),
    .B1(_00795_),
    .C1(_00797_),
    .Y(_01059_));
 sky130_fd_sc_hd__a211o_1 _07624_ (.A1(_00911_),
    .A2(_00913_),
    .B1(_01057_),
    .C1(_01059_),
    .X(_01060_));
 sky130_fd_sc_hd__o211ai_1 _07625_ (.A1(_01057_),
    .A2(_01059_),
    .B1(_00911_),
    .C1(_00913_),
    .Y(_01062_));
 sky130_fd_sc_hd__and3b_1 _07626_ (.A_N(_00915_),
    .B(_01060_),
    .C(_01062_),
    .X(_01063_));
 sky130_fd_sc_hd__a21boi_1 _07627_ (.A1(_01060_),
    .A2(_01062_),
    .B1_N(_00915_),
    .Y(_01064_));
 sky130_fd_sc_hd__nor2_2 _07628_ (.A(_01063_),
    .B(_01064_),
    .Y(_01065_));
 sky130_fd_sc_hd__nor2_1 _07629_ (.A(_00770_),
    .B(_00918_),
    .Y(_01066_));
 sky130_fd_sc_hd__nor2_1 _07630_ (.A(_00917_),
    .B(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__or3_1 _07631_ (.A(_00771_),
    .B(_00917_),
    .C(_00918_),
    .X(_01068_));
 sky130_fd_sc_hd__o21bai_2 _07632_ (.A1(_00777_),
    .A2(_01068_),
    .B1_N(_01067_),
    .Y(_01069_));
 sky130_fd_sc_hd__xor2_1 _07633_ (.A(_01065_),
    .B(_01069_),
    .X(net83));
 sky130_fd_sc_hd__a21o_1 _07634_ (.A1(_00782_),
    .A2(_00932_),
    .B1(_00931_),
    .X(_01070_));
 sky130_fd_sc_hd__a21oi_1 _07635_ (.A1(_00950_),
    .A2(_00959_),
    .B1(_00957_),
    .Y(_01072_));
 sky130_fd_sc_hd__nand2_1 _07636_ (.A(_00925_),
    .B(_00928_),
    .Y(_01073_));
 sky130_fd_sc_hd__o21ba_1 _07637_ (.A1(_00946_),
    .A2(_00948_),
    .B1_N(_00947_),
    .X(_01074_));
 sky130_fd_sc_hd__and4_1 _07638_ (.A(net26),
    .B(net23),
    .C(net49),
    .D(net50),
    .X(_01075_));
 sky130_fd_sc_hd__a22oi_1 _07639_ (.A1(net26),
    .A2(net49),
    .B1(net50),
    .B2(net23),
    .Y(_01076_));
 sky130_fd_sc_hd__nor2_1 _07640_ (.A(_01075_),
    .B(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__nand2_1 _07641_ (.A(net12),
    .B(net51),
    .Y(_01078_));
 sky130_fd_sc_hd__xnor2_1 _07642_ (.A(_01077_),
    .B(_01078_),
    .Y(_01079_));
 sky130_fd_sc_hd__nand2b_1 _07643_ (.A_N(_01074_),
    .B(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__xnor2_1 _07644_ (.A(_01074_),
    .B(_01079_),
    .Y(_01081_));
 sky130_fd_sc_hd__nand2_1 _07645_ (.A(_01073_),
    .B(_01081_),
    .Y(_01083_));
 sky130_fd_sc_hd__xor2_1 _07646_ (.A(_01073_),
    .B(_01081_),
    .X(_01084_));
 sky130_fd_sc_hd__and2b_1 _07647_ (.A_N(_01072_),
    .B(_01084_),
    .X(_01085_));
 sky130_fd_sc_hd__xnor2_1 _07648_ (.A(_01072_),
    .B(_01084_),
    .Y(_01086_));
 sky130_fd_sc_hd__and2_1 _07649_ (.A(_01070_),
    .B(_01086_),
    .X(_01087_));
 sky130_fd_sc_hd__xnor2_1 _07650_ (.A(_01070_),
    .B(_01086_),
    .Y(_01088_));
 sky130_fd_sc_hd__a21oi_1 _07651_ (.A1(_00784_),
    .A2(_00936_),
    .B1(_00935_),
    .Y(_01089_));
 sky130_fd_sc_hd__or2_1 _07652_ (.A(_01088_),
    .B(_01089_),
    .X(_01090_));
 sky130_fd_sc_hd__xnor2_1 _07653_ (.A(_01088_),
    .B(_01089_),
    .Y(_01091_));
 sky130_fd_sc_hd__nand2_1 _07654_ (.A(net1),
    .B(net52),
    .Y(_01092_));
 sky130_fd_sc_hd__or2_1 _07655_ (.A(_01091_),
    .B(_01092_),
    .X(_01094_));
 sky130_fd_sc_hd__xor2_1 _07656_ (.A(_01091_),
    .B(_01092_),
    .X(_01095_));
 sky130_fd_sc_hd__nor3_1 _07657_ (.A(_00979_),
    .B(_00981_),
    .C(_01095_),
    .Y(_01096_));
 sky130_fd_sc_hd__o21a_1 _07658_ (.A1(_00979_),
    .A2(_00981_),
    .B1(_01095_),
    .X(_01097_));
 sky130_fd_sc_hd__o21ai_2 _07659_ (.A1(_01096_),
    .A2(_01097_),
    .B1(_00938_),
    .Y(_01098_));
 sky130_fd_sc_hd__or3_2 _07660_ (.A(_00938_),
    .B(_01096_),
    .C(_01097_),
    .X(_01099_));
 sky130_fd_sc_hd__nand2_1 _07661_ (.A(net27),
    .B(net48),
    .Y(_01100_));
 sky130_fd_sc_hd__and4_1 _07662_ (.A(net28),
    .B(net29),
    .C(net46),
    .D(net47),
    .X(_01101_));
 sky130_fd_sc_hd__a22oi_1 _07663_ (.A1(net29),
    .A2(net46),
    .B1(net47),
    .B2(net28),
    .Y(_01102_));
 sky130_fd_sc_hd__nor2_1 _07664_ (.A(_01101_),
    .B(_01102_),
    .Y(_01103_));
 sky130_fd_sc_hd__xnor2_1 _07665_ (.A(_01100_),
    .B(_01103_),
    .Y(_01105_));
 sky130_fd_sc_hd__nand2_1 _07666_ (.A(net30),
    .B(net45),
    .Y(_01106_));
 sky130_fd_sc_hd__and4_1 _07667_ (.A(net31),
    .B(net32),
    .C(net42),
    .D(net43),
    .X(_01107_));
 sky130_fd_sc_hd__a22oi_1 _07668_ (.A1(net32),
    .A2(net42),
    .B1(net43),
    .B2(net31),
    .Y(_01108_));
 sky130_fd_sc_hd__nor2_1 _07669_ (.A(_01107_),
    .B(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__xnor2_1 _07670_ (.A(_01106_),
    .B(_01109_),
    .Y(_01110_));
 sky130_fd_sc_hd__nor2_1 _07671_ (.A(_00951_),
    .B(_00954_),
    .Y(_01111_));
 sky130_fd_sc_hd__and2b_1 _07672_ (.A_N(_01111_),
    .B(_01110_),
    .X(_01112_));
 sky130_fd_sc_hd__xnor2_1 _07673_ (.A(_01110_),
    .B(_01111_),
    .Y(_01113_));
 sky130_fd_sc_hd__and2_1 _07674_ (.A(_01105_),
    .B(_01113_),
    .X(_01114_));
 sky130_fd_sc_hd__nor2_1 _07675_ (.A(_01105_),
    .B(_01113_),
    .Y(_01116_));
 sky130_fd_sc_hd__or2_1 _07676_ (.A(_01114_),
    .B(_01116_),
    .X(_01117_));
 sky130_fd_sc_hd__a31o_1 _07677_ (.A1(net32),
    .A2(net41),
    .A3(_00966_),
    .B1(_00964_),
    .X(_01118_));
 sky130_fd_sc_hd__o21ba_1 _07678_ (.A1(_00983_),
    .A2(_00986_),
    .B1_N(_00985_),
    .X(_01119_));
 sky130_fd_sc_hd__nand2_1 _07679_ (.A(net2),
    .B(net41),
    .Y(_01120_));
 sky130_fd_sc_hd__and4_1 _07680_ (.A(net3),
    .B(net4),
    .C(net39),
    .D(net40),
    .X(_01121_));
 sky130_fd_sc_hd__a22oi_1 _07681_ (.A1(net4),
    .A2(net39),
    .B1(net40),
    .B2(net3),
    .Y(_01122_));
 sky130_fd_sc_hd__nor2_1 _07682_ (.A(_01121_),
    .B(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__xnor2_1 _07683_ (.A(_01120_),
    .B(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2b_1 _07684_ (.A_N(_01119_),
    .B(_01124_),
    .Y(_01125_));
 sky130_fd_sc_hd__xnor2_1 _07685_ (.A(_01119_),
    .B(_01124_),
    .Y(_01127_));
 sky130_fd_sc_hd__nand2_1 _07686_ (.A(_01118_),
    .B(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__xnor2_1 _07687_ (.A(_01118_),
    .B(_01127_),
    .Y(_01129_));
 sky130_fd_sc_hd__a21o_1 _07688_ (.A1(_00968_),
    .A2(_00970_),
    .B1(_01129_),
    .X(_01130_));
 sky130_fd_sc_hd__nand3_1 _07689_ (.A(_00968_),
    .B(_00970_),
    .C(_01129_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand3b_2 _07690_ (.A_N(_01117_),
    .B(_01130_),
    .C(_01131_),
    .Y(_01132_));
 sky130_fd_sc_hd__a21bo_1 _07691_ (.A1(_01130_),
    .A2(_01131_),
    .B1_N(_01117_),
    .X(_01133_));
 sky130_fd_sc_hd__o211a_1 _07692_ (.A1(_01000_),
    .A2(_01003_),
    .B1(_01132_),
    .C1(_01133_),
    .X(_01134_));
 sky130_fd_sc_hd__a211oi_1 _07693_ (.A1(_01132_),
    .A2(_01133_),
    .B1(_01000_),
    .C1(_01003_),
    .Y(_01135_));
 sky130_fd_sc_hd__a211oi_2 _07694_ (.A1(_00974_),
    .A2(_00977_),
    .B1(_01134_),
    .C1(_01135_),
    .Y(_01136_));
 sky130_fd_sc_hd__o211a_1 _07695_ (.A1(_01134_),
    .A2(_01135_),
    .B1(_00974_),
    .C1(_00977_),
    .X(_01138_));
 sky130_fd_sc_hd__nand2_1 _07696_ (.A(net5),
    .B(net38),
    .Y(_01139_));
 sky130_fd_sc_hd__and4_1 _07697_ (.A(net36),
    .B(net37),
    .C(net6),
    .D(net7),
    .X(_01140_));
 sky130_fd_sc_hd__a22oi_1 _07698_ (.A1(net37),
    .A2(net6),
    .B1(net7),
    .B2(net36),
    .Y(_01141_));
 sky130_fd_sc_hd__nor2_1 _07699_ (.A(_01140_),
    .B(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__xnor2_1 _07700_ (.A(_01139_),
    .B(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hd__and4_1 _07701_ (.A(net64),
    .B(net34),
    .C(net9),
    .D(net10),
    .X(_01144_));
 sky130_fd_sc_hd__a22oi_1 _07702_ (.A1(net34),
    .A2(net9),
    .B1(net10),
    .B2(net64),
    .Y(_01145_));
 sky130_fd_sc_hd__and4bb_1 _07703_ (.A_N(_01144_),
    .B_N(_01145_),
    .C(net35),
    .D(net8),
    .X(_01146_));
 sky130_fd_sc_hd__o2bb2a_1 _07704_ (.A1_N(net35),
    .A2_N(net8),
    .B1(_01144_),
    .B2(_01145_),
    .X(_01147_));
 sky130_fd_sc_hd__nor2_1 _07705_ (.A(_01146_),
    .B(_01147_),
    .Y(_01149_));
 sky130_fd_sc_hd__o21ba_1 _07706_ (.A1(_00989_),
    .A2(_00991_),
    .B1_N(_00990_),
    .X(_01150_));
 sky130_fd_sc_hd__and2b_1 _07707_ (.A_N(_01150_),
    .B(_01149_),
    .X(_01151_));
 sky130_fd_sc_hd__xnor2_1 _07708_ (.A(_01149_),
    .B(_01150_),
    .Y(_01152_));
 sky130_fd_sc_hd__and2_1 _07709_ (.A(_01143_),
    .B(_01152_),
    .X(_01153_));
 sky130_fd_sc_hd__xnor2_1 _07710_ (.A(_01143_),
    .B(_01152_),
    .Y(_01154_));
 sky130_fd_sc_hd__a21o_2 _07711_ (.A1(_01013_),
    .A2(_01015_),
    .B1(_01154_),
    .X(_01155_));
 sky130_fd_sc_hd__nand3_1 _07712_ (.A(_01013_),
    .B(_01015_),
    .C(_01154_),
    .Y(_01156_));
 sky130_fd_sc_hd__o211ai_4 _07713_ (.A1(_00996_),
    .A2(_00998_),
    .B1(_01155_),
    .C1(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__a211o_1 _07714_ (.A1(_01155_),
    .A2(_01156_),
    .B1(_00996_),
    .C1(_00998_),
    .X(_01158_));
 sky130_fd_sc_hd__o21ba_1 _07715_ (.A1(_01008_),
    .A2(_01010_),
    .B1_N(_01009_),
    .X(_01160_));
 sky130_fd_sc_hd__o21ba_1 _07716_ (.A1(_01018_),
    .A2(_01020_),
    .B1_N(_01019_),
    .X(_01161_));
 sky130_fd_sc_hd__nand2_1 _07717_ (.A(net63),
    .B(net11),
    .Y(_01162_));
 sky130_fd_sc_hd__and4_1 _07718_ (.A(net61),
    .B(net62),
    .C(net13),
    .D(net14),
    .X(_01163_));
 sky130_fd_sc_hd__a22oi_1 _07719_ (.A1(net62),
    .A2(net13),
    .B1(net14),
    .B2(net61),
    .Y(_01164_));
 sky130_fd_sc_hd__nor2_1 _07720_ (.A(_01163_),
    .B(_01164_),
    .Y(_01165_));
 sky130_fd_sc_hd__xnor2_1 _07721_ (.A(_01162_),
    .B(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__nand2b_1 _07722_ (.A_N(_01161_),
    .B(_01166_),
    .Y(_01167_));
 sky130_fd_sc_hd__xnor2_1 _07723_ (.A(_01161_),
    .B(_01166_),
    .Y(_01168_));
 sky130_fd_sc_hd__nand2b_1 _07724_ (.A_N(_01160_),
    .B(_01168_),
    .Y(_01169_));
 sky130_fd_sc_hd__xnor2_1 _07725_ (.A(_01160_),
    .B(_01168_),
    .Y(_01171_));
 sky130_fd_sc_hd__nand2_1 _07726_ (.A(net60),
    .B(net15),
    .Y(_01172_));
 sky130_fd_sc_hd__and4_1 _07727_ (.A(net58),
    .B(net59),
    .C(net16),
    .D(net17),
    .X(_01173_));
 sky130_fd_sc_hd__a22oi_1 _07728_ (.A1(net59),
    .A2(net16),
    .B1(net17),
    .B2(net58),
    .Y(_01174_));
 sky130_fd_sc_hd__nor2_1 _07729_ (.A(_01173_),
    .B(_01174_),
    .Y(_01175_));
 sky130_fd_sc_hd__xnor2_1 _07730_ (.A(_01172_),
    .B(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hd__and2_1 _07731_ (.A(net55),
    .B(net18),
    .X(_01177_));
 sky130_fd_sc_hd__nand4_1 _07732_ (.A(net33),
    .B(net44),
    .C(net19),
    .D(net20),
    .Y(_01178_));
 sky130_fd_sc_hd__a22o_1 _07733_ (.A1(net44),
    .A2(net19),
    .B1(net20),
    .B2(net33),
    .X(_01179_));
 sky130_fd_sc_hd__nand3_1 _07734_ (.A(_01177_),
    .B(_01178_),
    .C(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__a21o_1 _07735_ (.A1(_01178_),
    .A2(_01179_),
    .B1(_01177_),
    .X(_01182_));
 sky130_fd_sc_hd__o21bai_1 _07736_ (.A1(_01023_),
    .A2(_01025_),
    .B1_N(_01024_),
    .Y(_01183_));
 sky130_fd_sc_hd__nand3_1 _07737_ (.A(_01180_),
    .B(_01182_),
    .C(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__a21o_1 _07738_ (.A1(_01180_),
    .A2(_01182_),
    .B1(_01183_),
    .X(_01185_));
 sky130_fd_sc_hd__nand3_1 _07739_ (.A(_01176_),
    .B(_01184_),
    .C(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__a21o_1 _07740_ (.A1(_01184_),
    .A2(_01185_),
    .B1(_01176_),
    .X(_01187_));
 sky130_fd_sc_hd__a21bo_1 _07741_ (.A1(_01022_),
    .A2(_01031_),
    .B1_N(_01030_),
    .X(_01188_));
 sky130_fd_sc_hd__nand3_2 _07742_ (.A(_01186_),
    .B(_01187_),
    .C(_01188_),
    .Y(_01189_));
 sky130_fd_sc_hd__a21o_1 _07743_ (.A1(_01186_),
    .A2(_01187_),
    .B1(_01188_),
    .X(_01190_));
 sky130_fd_sc_hd__and3_1 _07744_ (.A(_01171_),
    .B(_01189_),
    .C(_01190_),
    .X(_01191_));
 sky130_fd_sc_hd__nand3_1 _07745_ (.A(_01171_),
    .B(_01189_),
    .C(_01190_),
    .Y(_01193_));
 sky130_fd_sc_hd__a21oi_2 _07746_ (.A1(_01189_),
    .A2(_01190_),
    .B1(_01171_),
    .Y(_01194_));
 sky130_fd_sc_hd__a211oi_2 _07747_ (.A1(_01035_),
    .A2(_01038_),
    .B1(_01191_),
    .C1(_01194_),
    .Y(_01195_));
 sky130_fd_sc_hd__a211o_1 _07748_ (.A1(_01035_),
    .A2(_01038_),
    .B1(_01191_),
    .C1(_01194_),
    .X(_01196_));
 sky130_fd_sc_hd__o211ai_2 _07749_ (.A1(_01191_),
    .A2(_01194_),
    .B1(_01035_),
    .C1(_01038_),
    .Y(_01197_));
 sky130_fd_sc_hd__and4_1 _07750_ (.A(_01157_),
    .B(_01158_),
    .C(_01196_),
    .D(_01197_),
    .X(_01198_));
 sky130_fd_sc_hd__a22oi_2 _07751_ (.A1(_01157_),
    .A2(_01158_),
    .B1(_01196_),
    .B2(_01197_),
    .Y(_01199_));
 sky130_fd_sc_hd__a211o_1 _07752_ (.A1(_01041_),
    .A2(_01043_),
    .B1(_01198_),
    .C1(_01199_),
    .X(_01200_));
 sky130_fd_sc_hd__o211ai_1 _07753_ (.A1(_01198_),
    .A2(_01199_),
    .B1(_01041_),
    .C1(_01043_),
    .Y(_01201_));
 sky130_fd_sc_hd__or4bb_4 _07754_ (.A(_01136_),
    .B(_01138_),
    .C_N(_01200_),
    .D_N(_01201_),
    .X(_01202_));
 sky130_fd_sc_hd__a2bb2o_1 _07755_ (.A1_N(_01136_),
    .A2_N(_01138_),
    .B1(_01200_),
    .B2(_01201_),
    .X(_01204_));
 sky130_fd_sc_hd__o211ai_4 _07756_ (.A1(_01045_),
    .A2(_01047_),
    .B1(_01202_),
    .C1(_01204_),
    .Y(_01205_));
 sky130_fd_sc_hd__a211o_1 _07757_ (.A1(_01202_),
    .A2(_01204_),
    .B1(_01045_),
    .C1(_01047_),
    .X(_01206_));
 sky130_fd_sc_hd__nand4_4 _07758_ (.A(_01098_),
    .B(_01099_),
    .C(_01205_),
    .D(_01206_),
    .Y(_01207_));
 sky130_fd_sc_hd__a22o_1 _07759_ (.A1(_01098_),
    .A2(_01099_),
    .B1(_01205_),
    .B2(_01206_),
    .X(_01208_));
 sky130_fd_sc_hd__o211a_2 _07760_ (.A1(_01049_),
    .A2(_01052_),
    .B1(_01207_),
    .C1(_01208_),
    .X(_01209_));
 sky130_fd_sc_hd__a211oi_2 _07761_ (.A1(_01207_),
    .A2(_01208_),
    .B1(_01049_),
    .C1(_01052_),
    .Y(_01210_));
 sky130_fd_sc_hd__a211oi_4 _07762_ (.A1(_00942_),
    .A2(_00944_),
    .B1(_01209_),
    .C1(_01210_),
    .Y(_01211_));
 sky130_fd_sc_hd__o211a_1 _07763_ (.A1(_01209_),
    .A2(_01210_),
    .B1(_00942_),
    .C1(_00944_),
    .X(_01212_));
 sky130_fd_sc_hd__a211oi_2 _07764_ (.A1(_01055_),
    .A2(_01058_),
    .B1(_01211_),
    .C1(_01212_),
    .Y(_01213_));
 sky130_fd_sc_hd__o211a_1 _07765_ (.A1(_01211_),
    .A2(_01212_),
    .B1(_01055_),
    .C1(_01058_),
    .X(_01215_));
 sky130_fd_sc_hd__o21a_1 _07766_ (.A1(_01213_),
    .A2(_01215_),
    .B1(_01060_),
    .X(_01216_));
 sky130_fd_sc_hd__nor3_1 _07767_ (.A(_01060_),
    .B(_01213_),
    .C(_01215_),
    .Y(_01217_));
 sky130_fd_sc_hd__nor2_1 _07768_ (.A(_01216_),
    .B(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__a21oi_1 _07769_ (.A1(_01065_),
    .A2(_01069_),
    .B1(_01063_),
    .Y(_01219_));
 sky130_fd_sc_hd__xnor2_1 _07770_ (.A(_01218_),
    .B(_01219_),
    .Y(net84));
 sky130_fd_sc_hd__o21ba_1 _07771_ (.A1(_01063_),
    .A2(_01217_),
    .B1_N(_01216_),
    .X(_01220_));
 sky130_fd_sc_hd__a31oi_4 _07772_ (.A1(_01065_),
    .A2(_01069_),
    .A3(_01218_),
    .B1(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__and2b_1 _07773_ (.A_N(_01097_),
    .B(_01099_),
    .X(_01222_));
 sky130_fd_sc_hd__a22o_1 _07774_ (.A1(net12),
    .A2(net52),
    .B1(net53),
    .B2(net1),
    .X(_01223_));
 sky130_fd_sc_hd__and4_1 _07775_ (.A(net12),
    .B(net1),
    .C(net52),
    .D(net53),
    .X(_01225_));
 sky130_fd_sc_hd__nand4_1 _07776_ (.A(net12),
    .B(net1),
    .C(net52),
    .D(net53),
    .Y(_01226_));
 sky130_fd_sc_hd__o21ba_1 _07777_ (.A1(_01076_),
    .A2(_01078_),
    .B1_N(_01075_),
    .X(_01227_));
 sky130_fd_sc_hd__o21ba_1 _07778_ (.A1(_01100_),
    .A2(_01102_),
    .B1_N(_01101_),
    .X(_01228_));
 sky130_fd_sc_hd__and4_1 _07779_ (.A(net27),
    .B(net26),
    .C(net49),
    .D(net50),
    .X(_01229_));
 sky130_fd_sc_hd__a22oi_1 _07780_ (.A1(net27),
    .A2(net49),
    .B1(net50),
    .B2(net26),
    .Y(_01230_));
 sky130_fd_sc_hd__nor2_1 _07781_ (.A(_01229_),
    .B(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__nand2_1 _07782_ (.A(net23),
    .B(net51),
    .Y(_01232_));
 sky130_fd_sc_hd__xnor2_1 _07783_ (.A(_01231_),
    .B(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__and2b_1 _07784_ (.A_N(_01228_),
    .B(_01233_),
    .X(_01234_));
 sky130_fd_sc_hd__xnor2_1 _07785_ (.A(_01228_),
    .B(_01233_),
    .Y(_01236_));
 sky130_fd_sc_hd__and2b_1 _07786_ (.A_N(_01227_),
    .B(_01236_),
    .X(_01237_));
 sky130_fd_sc_hd__xnor2_1 _07787_ (.A(_01227_),
    .B(_01236_),
    .Y(_01238_));
 sky130_fd_sc_hd__o21a_1 _07788_ (.A1(_01112_),
    .A2(_01114_),
    .B1(_01238_),
    .X(_01239_));
 sky130_fd_sc_hd__nor3_1 _07789_ (.A(_01112_),
    .B(_01114_),
    .C(_01238_),
    .Y(_01240_));
 sky130_fd_sc_hd__a211oi_1 _07790_ (.A1(_01080_),
    .A2(_01083_),
    .B1(_01239_),
    .C1(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__a211o_1 _07791_ (.A1(_01080_),
    .A2(_01083_),
    .B1(_01239_),
    .C1(_01240_),
    .X(_01242_));
 sky130_fd_sc_hd__o211ai_2 _07792_ (.A1(_01239_),
    .A2(_01240_),
    .B1(_01080_),
    .C1(_01083_),
    .Y(_01243_));
 sky130_fd_sc_hd__o211ai_4 _07793_ (.A1(_01085_),
    .A2(_01087_),
    .B1(_01242_),
    .C1(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hd__a211o_1 _07794_ (.A1(_01242_),
    .A2(_01243_),
    .B1(_01085_),
    .C1(_01087_),
    .X(_01245_));
 sky130_fd_sc_hd__nand4_2 _07795_ (.A(_01223_),
    .B(_01226_),
    .C(_01244_),
    .D(_01245_),
    .Y(_01247_));
 sky130_fd_sc_hd__a22o_1 _07796_ (.A1(_01223_),
    .A2(_01226_),
    .B1(_01244_),
    .B2(_01245_),
    .X(_01248_));
 sky130_fd_sc_hd__o211a_1 _07797_ (.A1(_01134_),
    .A2(_01136_),
    .B1(_01247_),
    .C1(_01248_),
    .X(_01249_));
 sky130_fd_sc_hd__inv_2 _07798_ (.A(_01249_),
    .Y(_01250_));
 sky130_fd_sc_hd__a211oi_1 _07799_ (.A1(_01247_),
    .A2(_01248_),
    .B1(_01134_),
    .C1(_01136_),
    .Y(_01251_));
 sky130_fd_sc_hd__a211o_1 _07800_ (.A1(_01090_),
    .A2(_01094_),
    .B1(_01249_),
    .C1(_01251_),
    .X(_01252_));
 sky130_fd_sc_hd__o211ai_1 _07801_ (.A1(_01249_),
    .A2(_01251_),
    .B1(_01090_),
    .C1(_01094_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand2_1 _07802_ (.A(net28),
    .B(net48),
    .Y(_01254_));
 sky130_fd_sc_hd__and4_1 _07803_ (.A(net29),
    .B(net30),
    .C(net46),
    .D(net47),
    .X(_01255_));
 sky130_fd_sc_hd__a22oi_1 _07804_ (.A1(net30),
    .A2(net46),
    .B1(net47),
    .B2(net29),
    .Y(_01256_));
 sky130_fd_sc_hd__nor2_1 _07805_ (.A(_01255_),
    .B(_01256_),
    .Y(_01258_));
 sky130_fd_sc_hd__xnor2_1 _07806_ (.A(_01254_),
    .B(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__nand2_1 _07807_ (.A(net31),
    .B(net45),
    .Y(_01260_));
 sky130_fd_sc_hd__and4_1 _07808_ (.A(net2),
    .B(net32),
    .C(net42),
    .D(net43),
    .X(_01261_));
 sky130_fd_sc_hd__a22oi_1 _07809_ (.A1(net2),
    .A2(net42),
    .B1(net43),
    .B2(net32),
    .Y(_01262_));
 sky130_fd_sc_hd__nor2_1 _07810_ (.A(_01261_),
    .B(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__xnor2_1 _07811_ (.A(_01260_),
    .B(_01263_),
    .Y(_01264_));
 sky130_fd_sc_hd__o21ba_1 _07812_ (.A1(_01106_),
    .A2(_01108_),
    .B1_N(_01107_),
    .X(_01265_));
 sky130_fd_sc_hd__and2b_1 _07813_ (.A_N(_01265_),
    .B(_01264_),
    .X(_01266_));
 sky130_fd_sc_hd__xnor2_1 _07814_ (.A(_01264_),
    .B(_01265_),
    .Y(_01267_));
 sky130_fd_sc_hd__and2_1 _07815_ (.A(_01259_),
    .B(_01267_),
    .X(_01269_));
 sky130_fd_sc_hd__nor2_1 _07816_ (.A(_01259_),
    .B(_01267_),
    .Y(_01270_));
 sky130_fd_sc_hd__or2_1 _07817_ (.A(_01269_),
    .B(_01270_),
    .X(_01271_));
 sky130_fd_sc_hd__a31o_1 _07818_ (.A1(net2),
    .A2(net41),
    .A3(_01123_),
    .B1(_01121_),
    .X(_01272_));
 sky130_fd_sc_hd__o21ba_1 _07819_ (.A1(_01139_),
    .A2(_01141_),
    .B1_N(_01140_),
    .X(_01273_));
 sky130_fd_sc_hd__a22oi_1 _07820_ (.A1(net5),
    .A2(net39),
    .B1(net40),
    .B2(net4),
    .Y(_01274_));
 sky130_fd_sc_hd__and4_1 _07821_ (.A(net4),
    .B(net5),
    .C(net39),
    .D(net40),
    .X(_01275_));
 sky130_fd_sc_hd__nor2_1 _07822_ (.A(_01274_),
    .B(_01275_),
    .Y(_01276_));
 sky130_fd_sc_hd__nand2_1 _07823_ (.A(net3),
    .B(net41),
    .Y(_01277_));
 sky130_fd_sc_hd__xnor2_1 _07824_ (.A(_01276_),
    .B(_01277_),
    .Y(_01278_));
 sky130_fd_sc_hd__nand2b_1 _07825_ (.A_N(_01273_),
    .B(_01278_),
    .Y(_01280_));
 sky130_fd_sc_hd__xnor2_1 _07826_ (.A(_01273_),
    .B(_01278_),
    .Y(_01281_));
 sky130_fd_sc_hd__nand2_1 _07827_ (.A(_01272_),
    .B(_01281_),
    .Y(_01282_));
 sky130_fd_sc_hd__xnor2_1 _07828_ (.A(_01272_),
    .B(_01281_),
    .Y(_01283_));
 sky130_fd_sc_hd__a21oi_1 _07829_ (.A1(_01125_),
    .A2(_01128_),
    .B1(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__and3_1 _07830_ (.A(_01125_),
    .B(_01128_),
    .C(_01283_),
    .X(_01285_));
 sky130_fd_sc_hd__nor3_1 _07831_ (.A(_01271_),
    .B(_01284_),
    .C(_01285_),
    .Y(_01286_));
 sky130_fd_sc_hd__o21a_1 _07832_ (.A1(_01284_),
    .A2(_01285_),
    .B1(_01271_),
    .X(_01287_));
 sky130_fd_sc_hd__a211oi_2 _07833_ (.A1(_01155_),
    .A2(_01157_),
    .B1(_01286_),
    .C1(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__o211a_1 _07834_ (.A1(_01286_),
    .A2(_01287_),
    .B1(_01155_),
    .C1(_01157_),
    .X(_01289_));
 sky130_fd_sc_hd__a211oi_2 _07835_ (.A1(_01130_),
    .A2(_01132_),
    .B1(_01288_),
    .C1(_01289_),
    .Y(_01291_));
 sky130_fd_sc_hd__o211a_1 _07836_ (.A1(_01288_),
    .A2(_01289_),
    .B1(_01130_),
    .C1(_01132_),
    .X(_01292_));
 sky130_fd_sc_hd__nand2_1 _07837_ (.A(net6),
    .B(net38),
    .Y(_01293_));
 sky130_fd_sc_hd__and4_1 _07838_ (.A(net36),
    .B(net37),
    .C(net7),
    .D(net8),
    .X(_01294_));
 sky130_fd_sc_hd__a22oi_1 _07839_ (.A1(net37),
    .A2(net7),
    .B1(net8),
    .B2(net36),
    .Y(_01295_));
 sky130_fd_sc_hd__nor2_1 _07840_ (.A(_01294_),
    .B(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hd__xnor2_1 _07841_ (.A(_01293_),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_1 _07842_ (.A(net35),
    .B(net9),
    .Y(_01298_));
 sky130_fd_sc_hd__and4_1 _07843_ (.A(net64),
    .B(net34),
    .C(net10),
    .D(net11),
    .X(_01299_));
 sky130_fd_sc_hd__a22oi_1 _07844_ (.A1(net34),
    .A2(net10),
    .B1(net11),
    .B2(net64),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_1 _07845_ (.A(_01299_),
    .B(_01300_),
    .Y(_01302_));
 sky130_fd_sc_hd__xnor2_1 _07846_ (.A(_01298_),
    .B(_01302_),
    .Y(_01303_));
 sky130_fd_sc_hd__nor2_1 _07847_ (.A(_01144_),
    .B(_01146_),
    .Y(_01304_));
 sky130_fd_sc_hd__and2b_1 _07848_ (.A_N(_01304_),
    .B(_01303_),
    .X(_01305_));
 sky130_fd_sc_hd__xnor2_1 _07849_ (.A(_01303_),
    .B(_01304_),
    .Y(_01306_));
 sky130_fd_sc_hd__and2_1 _07850_ (.A(_01297_),
    .B(_01306_),
    .X(_01307_));
 sky130_fd_sc_hd__xnor2_1 _07851_ (.A(_01297_),
    .B(_01306_),
    .Y(_01308_));
 sky130_fd_sc_hd__a21oi_1 _07852_ (.A1(_01167_),
    .A2(_01169_),
    .B1(_01308_),
    .Y(_01309_));
 sky130_fd_sc_hd__a21o_1 _07853_ (.A1(_01167_),
    .A2(_01169_),
    .B1(_01308_),
    .X(_01310_));
 sky130_fd_sc_hd__nand3_1 _07854_ (.A(_01167_),
    .B(_01169_),
    .C(_01308_),
    .Y(_01311_));
 sky130_fd_sc_hd__o211a_1 _07855_ (.A1(_01151_),
    .A2(_01153_),
    .B1(_01310_),
    .C1(_01311_),
    .X(_01313_));
 sky130_fd_sc_hd__a211oi_1 _07856_ (.A1(_01310_),
    .A2(_01311_),
    .B1(_01151_),
    .C1(_01153_),
    .Y(_01314_));
 sky130_fd_sc_hd__o21ba_1 _07857_ (.A1(_01162_),
    .A2(_01164_),
    .B1_N(_01163_),
    .X(_01315_));
 sky130_fd_sc_hd__o21ba_1 _07858_ (.A1(_01172_),
    .A2(_01174_),
    .B1_N(_01173_),
    .X(_01316_));
 sky130_fd_sc_hd__nand2_1 _07859_ (.A(net63),
    .B(net13),
    .Y(_01317_));
 sky130_fd_sc_hd__and4_1 _07860_ (.A(net61),
    .B(net62),
    .C(net14),
    .D(net15),
    .X(_01318_));
 sky130_fd_sc_hd__a22oi_1 _07861_ (.A1(net62),
    .A2(net14),
    .B1(net15),
    .B2(net61),
    .Y(_01319_));
 sky130_fd_sc_hd__nor2_1 _07862_ (.A(_01318_),
    .B(_01319_),
    .Y(_01320_));
 sky130_fd_sc_hd__xnor2_1 _07863_ (.A(_01317_),
    .B(_01320_),
    .Y(_01321_));
 sky130_fd_sc_hd__nand2b_1 _07864_ (.A_N(_01316_),
    .B(_01321_),
    .Y(_01322_));
 sky130_fd_sc_hd__xnor2_1 _07865_ (.A(_01316_),
    .B(_01321_),
    .Y(_01323_));
 sky130_fd_sc_hd__nand2b_1 _07866_ (.A_N(_01315_),
    .B(_01323_),
    .Y(_01324_));
 sky130_fd_sc_hd__xnor2_1 _07867_ (.A(_01315_),
    .B(_01323_),
    .Y(_01325_));
 sky130_fd_sc_hd__nand2_1 _07868_ (.A(net60),
    .B(net16),
    .Y(_01326_));
 sky130_fd_sc_hd__and4_1 _07869_ (.A(net58),
    .B(net59),
    .C(net17),
    .D(net18),
    .X(_01327_));
 sky130_fd_sc_hd__a22oi_1 _07870_ (.A1(net59),
    .A2(net17),
    .B1(net18),
    .B2(net58),
    .Y(_01328_));
 sky130_fd_sc_hd__nor2_1 _07871_ (.A(_01327_),
    .B(_01328_),
    .Y(_01329_));
 sky130_fd_sc_hd__xnor2_1 _07872_ (.A(_01326_),
    .B(_01329_),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_1 _07873_ (.A(net55),
    .B(net19),
    .Y(_01331_));
 sky130_fd_sc_hd__and4_1 _07874_ (.A(net33),
    .B(net44),
    .C(net20),
    .D(net21),
    .X(_01332_));
 sky130_fd_sc_hd__a22oi_2 _07875_ (.A1(net44),
    .A2(net20),
    .B1(net21),
    .B2(net33),
    .Y(_01334_));
 sky130_fd_sc_hd__or3_1 _07876_ (.A(_01331_),
    .B(_01332_),
    .C(_01334_),
    .X(_01335_));
 sky130_fd_sc_hd__o21ai_1 _07877_ (.A1(_01332_),
    .A2(_01334_),
    .B1(_01331_),
    .Y(_01336_));
 sky130_fd_sc_hd__a21bo_1 _07878_ (.A1(_01177_),
    .A2(_01179_),
    .B1_N(_01178_),
    .X(_01337_));
 sky130_fd_sc_hd__nand3_1 _07879_ (.A(_01335_),
    .B(_01336_),
    .C(_01337_),
    .Y(_01338_));
 sky130_fd_sc_hd__a21o_1 _07880_ (.A1(_01335_),
    .A2(_01336_),
    .B1(_01337_),
    .X(_01339_));
 sky130_fd_sc_hd__nand3_1 _07881_ (.A(_01330_),
    .B(_01338_),
    .C(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__a21o_1 _07882_ (.A1(_01338_),
    .A2(_01339_),
    .B1(_01330_),
    .X(_01341_));
 sky130_fd_sc_hd__a21bo_1 _07883_ (.A1(_01176_),
    .A2(_01185_),
    .B1_N(_01184_),
    .X(_01342_));
 sky130_fd_sc_hd__nand3_2 _07884_ (.A(_01340_),
    .B(_01341_),
    .C(_01342_),
    .Y(_01343_));
 sky130_fd_sc_hd__a21o_1 _07885_ (.A1(_01340_),
    .A2(_01341_),
    .B1(_01342_),
    .X(_01345_));
 sky130_fd_sc_hd__and3_1 _07886_ (.A(_01325_),
    .B(_01343_),
    .C(_01345_),
    .X(_01346_));
 sky130_fd_sc_hd__nand3_1 _07887_ (.A(_01325_),
    .B(_01343_),
    .C(_01345_),
    .Y(_01347_));
 sky130_fd_sc_hd__a21oi_1 _07888_ (.A1(_01343_),
    .A2(_01345_),
    .B1(_01325_),
    .Y(_01348_));
 sky130_fd_sc_hd__a211o_1 _07889_ (.A1(_01189_),
    .A2(_01193_),
    .B1(_01346_),
    .C1(_01348_),
    .X(_01349_));
 sky130_fd_sc_hd__o211ai_1 _07890_ (.A1(_01346_),
    .A2(_01348_),
    .B1(_01189_),
    .C1(_01193_),
    .Y(_01350_));
 sky130_fd_sc_hd__or4bb_2 _07891_ (.A(_01313_),
    .B(_01314_),
    .C_N(_01349_),
    .D_N(_01350_),
    .X(_01351_));
 sky130_fd_sc_hd__a2bb2o_1 _07892_ (.A1_N(_01313_),
    .A2_N(_01314_),
    .B1(_01349_),
    .B2(_01350_),
    .X(_01352_));
 sky130_fd_sc_hd__o211a_1 _07893_ (.A1(_01195_),
    .A2(_01198_),
    .B1(_01351_),
    .C1(_01352_),
    .X(_01353_));
 sky130_fd_sc_hd__a211oi_2 _07894_ (.A1(_01351_),
    .A2(_01352_),
    .B1(_01195_),
    .C1(_01198_),
    .Y(_01354_));
 sky130_fd_sc_hd__nor4_2 _07895_ (.A(_01291_),
    .B(_01292_),
    .C(_01353_),
    .D(_01354_),
    .Y(_01356_));
 sky130_fd_sc_hd__o22a_1 _07896_ (.A1(_01291_),
    .A2(_01292_),
    .B1(_01353_),
    .B2(_01354_),
    .X(_01357_));
 sky130_fd_sc_hd__a211oi_1 _07897_ (.A1(_01200_),
    .A2(_01202_),
    .B1(_01356_),
    .C1(_01357_),
    .Y(_01358_));
 sky130_fd_sc_hd__a211o_1 _07898_ (.A1(_01200_),
    .A2(_01202_),
    .B1(_01356_),
    .C1(_01357_),
    .X(_01359_));
 sky130_fd_sc_hd__o211ai_1 _07899_ (.A1(_01356_),
    .A2(_01357_),
    .B1(_01200_),
    .C1(_01202_),
    .Y(_01360_));
 sky130_fd_sc_hd__and4_1 _07900_ (.A(_01252_),
    .B(_01253_),
    .C(_01359_),
    .D(_01360_),
    .X(_01361_));
 sky130_fd_sc_hd__a22oi_2 _07901_ (.A1(_01252_),
    .A2(_01253_),
    .B1(_01359_),
    .B2(_01360_),
    .Y(_01362_));
 sky130_fd_sc_hd__a211oi_1 _07902_ (.A1(_01205_),
    .A2(_01207_),
    .B1(_01361_),
    .C1(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hd__a211o_1 _07903_ (.A1(_01205_),
    .A2(_01207_),
    .B1(_01361_),
    .C1(_01362_),
    .X(_01364_));
 sky130_fd_sc_hd__o211a_1 _07904_ (.A1(_01361_),
    .A2(_01362_),
    .B1(_01205_),
    .C1(_01207_),
    .X(_01365_));
 sky130_fd_sc_hd__or3_2 _07905_ (.A(_01222_),
    .B(_01363_),
    .C(_01365_),
    .X(_01367_));
 sky130_fd_sc_hd__o21ai_1 _07906_ (.A1(_01363_),
    .A2(_01365_),
    .B1(_01222_),
    .Y(_01368_));
 sky130_fd_sc_hd__o211a_1 _07907_ (.A1(_01209_),
    .A2(_01211_),
    .B1(_01367_),
    .C1(_01368_),
    .X(_01369_));
 sky130_fd_sc_hd__o211ai_1 _07908_ (.A1(_01209_),
    .A2(_01211_),
    .B1(_01367_),
    .C1(_01368_),
    .Y(_01370_));
 sky130_fd_sc_hd__a211o_1 _07909_ (.A1(_01367_),
    .A2(_01368_),
    .B1(_01209_),
    .C1(_01211_),
    .X(_01371_));
 sky130_fd_sc_hd__and3_1 _07910_ (.A(_01213_),
    .B(_01370_),
    .C(_01371_),
    .X(_01372_));
 sky130_fd_sc_hd__a21oi_1 _07911_ (.A1(_01370_),
    .A2(_01371_),
    .B1(_01213_),
    .Y(_01373_));
 sky130_fd_sc_hd__nor2_1 _07912_ (.A(_01372_),
    .B(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__xnor2_1 _07913_ (.A(_01221_),
    .B(_01374_),
    .Y(net85));
 sky130_fd_sc_hd__and4_1 _07914_ (.A(net23),
    .B(net12),
    .C(net52),
    .D(net53),
    .X(_01375_));
 sky130_fd_sc_hd__a22oi_1 _07915_ (.A1(net23),
    .A2(net52),
    .B1(net53),
    .B2(net12),
    .Y(_01377_));
 sky130_fd_sc_hd__nor2_1 _07916_ (.A(_01375_),
    .B(_01377_),
    .Y(_01378_));
 sky130_fd_sc_hd__nand2_1 _07917_ (.A(net1),
    .B(net54),
    .Y(_01379_));
 sky130_fd_sc_hd__xnor2_1 _07918_ (.A(_01378_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__nand2_1 _07919_ (.A(_01225_),
    .B(_01380_),
    .Y(_01381_));
 sky130_fd_sc_hd__or2_1 _07920_ (.A(_01225_),
    .B(_01380_),
    .X(_01382_));
 sky130_fd_sc_hd__nand2_1 _07921_ (.A(_01381_),
    .B(_01382_),
    .Y(_01383_));
 sky130_fd_sc_hd__o21ba_1 _07922_ (.A1(_01230_),
    .A2(_01232_),
    .B1_N(_01229_),
    .X(_01384_));
 sky130_fd_sc_hd__o21ba_1 _07923_ (.A1(_01254_),
    .A2(_01256_),
    .B1_N(_01255_),
    .X(_01385_));
 sky130_fd_sc_hd__and4_1 _07924_ (.A(net28),
    .B(net27),
    .C(net49),
    .D(net50),
    .X(_01386_));
 sky130_fd_sc_hd__a22oi_1 _07925_ (.A1(net28),
    .A2(net49),
    .B1(net50),
    .B2(net27),
    .Y(_01388_));
 sky130_fd_sc_hd__o2bb2a_1 _07926_ (.A1_N(net26),
    .A2_N(net51),
    .B1(_01386_),
    .B2(_01388_),
    .X(_01389_));
 sky130_fd_sc_hd__and4bb_1 _07927_ (.A_N(_01386_),
    .B_N(_01388_),
    .C(net26),
    .D(net51),
    .X(_01390_));
 sky130_fd_sc_hd__nor2_1 _07928_ (.A(_01389_),
    .B(_01390_),
    .Y(_01391_));
 sky130_fd_sc_hd__or3_1 _07929_ (.A(_01385_),
    .B(_01389_),
    .C(_01390_),
    .X(_01392_));
 sky130_fd_sc_hd__xnor2_1 _07930_ (.A(_01385_),
    .B(_01391_),
    .Y(_01393_));
 sky130_fd_sc_hd__nand2b_1 _07931_ (.A_N(_01384_),
    .B(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__xnor2_1 _07932_ (.A(_01384_),
    .B(_01393_),
    .Y(_01395_));
 sky130_fd_sc_hd__o21ai_4 _07933_ (.A1(_01266_),
    .A2(_01269_),
    .B1(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__or3_2 _07934_ (.A(_01266_),
    .B(_01269_),
    .C(_01395_),
    .X(_01397_));
 sky130_fd_sc_hd__o211ai_4 _07935_ (.A1(_01234_),
    .A2(_01237_),
    .B1(_01396_),
    .C1(_01397_),
    .Y(_01399_));
 sky130_fd_sc_hd__a211o_1 _07936_ (.A1(_01396_),
    .A2(_01397_),
    .B1(_01234_),
    .C1(_01237_),
    .X(_01400_));
 sky130_fd_sc_hd__o211a_1 _07937_ (.A1(_01239_),
    .A2(_01241_),
    .B1(_01399_),
    .C1(_01400_),
    .X(_01401_));
 sky130_fd_sc_hd__a211oi_1 _07938_ (.A1(_01399_),
    .A2(_01400_),
    .B1(_01239_),
    .C1(_01241_),
    .Y(_01402_));
 sky130_fd_sc_hd__or3_1 _07939_ (.A(_01383_),
    .B(_01401_),
    .C(_01402_),
    .X(_01403_));
 sky130_fd_sc_hd__o21ai_1 _07940_ (.A1(_01401_),
    .A2(_01402_),
    .B1(_01383_),
    .Y(_01404_));
 sky130_fd_sc_hd__o211a_1 _07941_ (.A1(_01288_),
    .A2(_01291_),
    .B1(_01403_),
    .C1(_01404_),
    .X(_01405_));
 sky130_fd_sc_hd__a211oi_1 _07942_ (.A1(_01403_),
    .A2(_01404_),
    .B1(_01288_),
    .C1(_01291_),
    .Y(_01406_));
 sky130_fd_sc_hd__a211oi_2 _07943_ (.A1(_01244_),
    .A2(_01247_),
    .B1(_01405_),
    .C1(_01406_),
    .Y(_01407_));
 sky130_fd_sc_hd__o211a_1 _07944_ (.A1(_01405_),
    .A2(_01406_),
    .B1(_01244_),
    .C1(_01247_),
    .X(_01408_));
 sky130_fd_sc_hd__nor2_1 _07945_ (.A(_01284_),
    .B(_01286_),
    .Y(_01410_));
 sky130_fd_sc_hd__and4_1 _07946_ (.A(net30),
    .B(net31),
    .C(net46),
    .D(net47),
    .X(_01411_));
 sky130_fd_sc_hd__a22oi_1 _07947_ (.A1(net31),
    .A2(net46),
    .B1(net47),
    .B2(net30),
    .Y(_01412_));
 sky130_fd_sc_hd__o2bb2a_1 _07948_ (.A1_N(net29),
    .A2_N(net48),
    .B1(_01411_),
    .B2(_01412_),
    .X(_01413_));
 sky130_fd_sc_hd__and4bb_1 _07949_ (.A_N(_01411_),
    .B_N(_01412_),
    .C(net29),
    .D(net48),
    .X(_01414_));
 sky130_fd_sc_hd__nor2_1 _07950_ (.A(_01413_),
    .B(_01414_),
    .Y(_01415_));
 sky130_fd_sc_hd__nand2_1 _07951_ (.A(net32),
    .B(net45),
    .Y(_01416_));
 sky130_fd_sc_hd__and4_1 _07952_ (.A(net2),
    .B(net3),
    .C(net42),
    .D(net43),
    .X(_01417_));
 sky130_fd_sc_hd__a22oi_1 _07953_ (.A1(net3),
    .A2(net42),
    .B1(net43),
    .B2(net2),
    .Y(_01418_));
 sky130_fd_sc_hd__nor2_1 _07954_ (.A(_01417_),
    .B(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__xnor2_1 _07955_ (.A(_01416_),
    .B(_01419_),
    .Y(_01421_));
 sky130_fd_sc_hd__o21ba_1 _07956_ (.A1(_01260_),
    .A2(_01262_),
    .B1_N(_01261_),
    .X(_01422_));
 sky130_fd_sc_hd__and2b_1 _07957_ (.A_N(_01422_),
    .B(_01421_),
    .X(_01423_));
 sky130_fd_sc_hd__xnor2_1 _07958_ (.A(_01421_),
    .B(_01422_),
    .Y(_01424_));
 sky130_fd_sc_hd__and2_1 _07959_ (.A(_01415_),
    .B(_01424_),
    .X(_01425_));
 sky130_fd_sc_hd__nor2_1 _07960_ (.A(_01415_),
    .B(_01424_),
    .Y(_01426_));
 sky130_fd_sc_hd__or2_1 _07961_ (.A(_01425_),
    .B(_01426_),
    .X(_01427_));
 sky130_fd_sc_hd__a31o_1 _07962_ (.A1(net3),
    .A2(net41),
    .A3(_01276_),
    .B1(_01275_),
    .X(_01428_));
 sky130_fd_sc_hd__o21ba_1 _07963_ (.A1(_01293_),
    .A2(_01295_),
    .B1_N(_01294_),
    .X(_01429_));
 sky130_fd_sc_hd__and4_1 _07964_ (.A(net5),
    .B(net6),
    .C(net39),
    .D(net40),
    .X(_01430_));
 sky130_fd_sc_hd__a22oi_1 _07965_ (.A1(net6),
    .A2(net39),
    .B1(net40),
    .B2(net5),
    .Y(_01432_));
 sky130_fd_sc_hd__nor2_1 _07966_ (.A(_01430_),
    .B(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_1 _07967_ (.A(net4),
    .B(net41),
    .Y(_01434_));
 sky130_fd_sc_hd__xnor2_1 _07968_ (.A(_01433_),
    .B(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2b_1 _07969_ (.A_N(_01429_),
    .B(_01435_),
    .Y(_01436_));
 sky130_fd_sc_hd__xnor2_1 _07970_ (.A(_01429_),
    .B(_01435_),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_1 _07971_ (.A(_01428_),
    .B(_01437_),
    .Y(_01438_));
 sky130_fd_sc_hd__xnor2_1 _07972_ (.A(_01428_),
    .B(_01437_),
    .Y(_01439_));
 sky130_fd_sc_hd__a21o_1 _07973_ (.A1(_01280_),
    .A2(_01282_),
    .B1(_01439_),
    .X(_01440_));
 sky130_fd_sc_hd__nand3_1 _07974_ (.A(_01280_),
    .B(_01282_),
    .C(_01439_),
    .Y(_01441_));
 sky130_fd_sc_hd__nand3b_2 _07975_ (.A_N(_01427_),
    .B(_01440_),
    .C(_01441_),
    .Y(_01443_));
 sky130_fd_sc_hd__a21bo_1 _07976_ (.A1(_01440_),
    .A2(_01441_),
    .B1_N(_01427_),
    .X(_01444_));
 sky130_fd_sc_hd__o211a_2 _07977_ (.A1(_01309_),
    .A2(_01313_),
    .B1(_01443_),
    .C1(_01444_),
    .X(_01445_));
 sky130_fd_sc_hd__a211oi_1 _07978_ (.A1(_01443_),
    .A2(_01444_),
    .B1(_01309_),
    .C1(_01313_),
    .Y(_01446_));
 sky130_fd_sc_hd__nor3_2 _07979_ (.A(_01410_),
    .B(_01445_),
    .C(_01446_),
    .Y(_01447_));
 sky130_fd_sc_hd__o21a_1 _07980_ (.A1(_01445_),
    .A2(_01446_),
    .B1(_01410_),
    .X(_01448_));
 sky130_fd_sc_hd__nand2_1 _07981_ (.A(net38),
    .B(net7),
    .Y(_01449_));
 sky130_fd_sc_hd__and4_1 _07982_ (.A(net36),
    .B(net37),
    .C(net8),
    .D(net9),
    .X(_01450_));
 sky130_fd_sc_hd__a22oi_1 _07983_ (.A1(net37),
    .A2(net8),
    .B1(net9),
    .B2(net36),
    .Y(_01451_));
 sky130_fd_sc_hd__nor2_1 _07984_ (.A(_01450_),
    .B(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__xnor2_1 _07985_ (.A(_01449_),
    .B(_01452_),
    .Y(_01454_));
 sky130_fd_sc_hd__nand2_1 _07986_ (.A(net35),
    .B(net10),
    .Y(_01455_));
 sky130_fd_sc_hd__and4_1 _07987_ (.A(net64),
    .B(net34),
    .C(net11),
    .D(net13),
    .X(_01456_));
 sky130_fd_sc_hd__a22o_1 _07988_ (.A1(net34),
    .A2(net11),
    .B1(net13),
    .B2(net64),
    .X(_01457_));
 sky130_fd_sc_hd__and2b_1 _07989_ (.A_N(_01456_),
    .B(_01457_),
    .X(_01458_));
 sky130_fd_sc_hd__xnor2_1 _07990_ (.A(_01455_),
    .B(_01458_),
    .Y(_01459_));
 sky130_fd_sc_hd__o21ba_1 _07991_ (.A1(_01298_),
    .A2(_01300_),
    .B1_N(_01299_),
    .X(_01460_));
 sky130_fd_sc_hd__and2b_1 _07992_ (.A_N(_01460_),
    .B(_01459_),
    .X(_01461_));
 sky130_fd_sc_hd__xnor2_1 _07993_ (.A(_01459_),
    .B(_01460_),
    .Y(_01462_));
 sky130_fd_sc_hd__and2_1 _07994_ (.A(_01454_),
    .B(_01462_),
    .X(_01463_));
 sky130_fd_sc_hd__xnor2_1 _07995_ (.A(_01454_),
    .B(_01462_),
    .Y(_01465_));
 sky130_fd_sc_hd__a21o_2 _07996_ (.A1(_01322_),
    .A2(_01324_),
    .B1(_01465_),
    .X(_01466_));
 sky130_fd_sc_hd__nand3_1 _07997_ (.A(_01322_),
    .B(_01324_),
    .C(_01465_),
    .Y(_01467_));
 sky130_fd_sc_hd__o211ai_4 _07998_ (.A1(_01305_),
    .A2(_01307_),
    .B1(_01466_),
    .C1(_01467_),
    .Y(_01468_));
 sky130_fd_sc_hd__a211o_1 _07999_ (.A1(_01466_),
    .A2(_01467_),
    .B1(_01305_),
    .C1(_01307_),
    .X(_01469_));
 sky130_fd_sc_hd__a31o_1 _08000_ (.A1(net63),
    .A2(net13),
    .A3(_01320_),
    .B1(_01318_),
    .X(_01470_));
 sky130_fd_sc_hd__o21bai_1 _08001_ (.A1(_01326_),
    .A2(_01328_),
    .B1_N(_01327_),
    .Y(_01471_));
 sky130_fd_sc_hd__nand2_1 _08002_ (.A(net63),
    .B(net14),
    .Y(_01472_));
 sky130_fd_sc_hd__nand4_1 _08003_ (.A(net61),
    .B(net62),
    .C(net15),
    .D(net16),
    .Y(_01473_));
 sky130_fd_sc_hd__a22o_1 _08004_ (.A1(net62),
    .A2(net15),
    .B1(net16),
    .B2(net61),
    .X(_01474_));
 sky130_fd_sc_hd__nand3b_1 _08005_ (.A_N(_01472_),
    .B(_01473_),
    .C(_01474_),
    .Y(_01476_));
 sky130_fd_sc_hd__a21bo_1 _08006_ (.A1(_01473_),
    .A2(_01474_),
    .B1_N(_01472_),
    .X(_01477_));
 sky130_fd_sc_hd__and3_1 _08007_ (.A(_01471_),
    .B(_01476_),
    .C(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__a21o_1 _08008_ (.A1(_01476_),
    .A2(_01477_),
    .B1(_01471_),
    .X(_01479_));
 sky130_fd_sc_hd__and2b_1 _08009_ (.A_N(_01478_),
    .B(_01479_),
    .X(_01480_));
 sky130_fd_sc_hd__xor2_1 _08010_ (.A(_01470_),
    .B(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__nand2_1 _08011_ (.A(net60),
    .B(net17),
    .Y(_01482_));
 sky130_fd_sc_hd__and4_1 _08012_ (.A(net58),
    .B(net59),
    .C(net18),
    .D(net19),
    .X(_01483_));
 sky130_fd_sc_hd__a22oi_1 _08013_ (.A1(net59),
    .A2(net18),
    .B1(net19),
    .B2(net58),
    .Y(_01484_));
 sky130_fd_sc_hd__nor2_1 _08014_ (.A(_01483_),
    .B(_01484_),
    .Y(_01485_));
 sky130_fd_sc_hd__xnor2_1 _08015_ (.A(_01482_),
    .B(_01485_),
    .Y(_01487_));
 sky130_fd_sc_hd__and2_1 _08016_ (.A(net55),
    .B(net20),
    .X(_01488_));
 sky130_fd_sc_hd__nand4_1 _08017_ (.A(net33),
    .B(net44),
    .C(net21),
    .D(net22),
    .Y(_01489_));
 sky130_fd_sc_hd__a22o_1 _08018_ (.A1(net44),
    .A2(net21),
    .B1(net22),
    .B2(net33),
    .X(_01490_));
 sky130_fd_sc_hd__nand3_1 _08019_ (.A(_01488_),
    .B(_01489_),
    .C(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__a21o_1 _08020_ (.A1(_01489_),
    .A2(_01490_),
    .B1(_01488_),
    .X(_01492_));
 sky130_fd_sc_hd__o21bai_1 _08021_ (.A1(_01331_),
    .A2(_01334_),
    .B1_N(_01332_),
    .Y(_01493_));
 sky130_fd_sc_hd__nand3_1 _08022_ (.A(_01491_),
    .B(_01492_),
    .C(_01493_),
    .Y(_01494_));
 sky130_fd_sc_hd__a21o_1 _08023_ (.A1(_01491_),
    .A2(_01492_),
    .B1(_01493_),
    .X(_01495_));
 sky130_fd_sc_hd__nand3_1 _08024_ (.A(_01487_),
    .B(_01494_),
    .C(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__a21o_1 _08025_ (.A1(_01494_),
    .A2(_01495_),
    .B1(_01487_),
    .X(_01498_));
 sky130_fd_sc_hd__a21bo_1 _08026_ (.A1(_01330_),
    .A2(_01339_),
    .B1_N(_01338_),
    .X(_01499_));
 sky130_fd_sc_hd__nand3_2 _08027_ (.A(_01496_),
    .B(_01498_),
    .C(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__a21o_1 _08028_ (.A1(_01496_),
    .A2(_01498_),
    .B1(_01499_),
    .X(_01501_));
 sky130_fd_sc_hd__and3_1 _08029_ (.A(_01481_),
    .B(_01500_),
    .C(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__nand3_1 _08030_ (.A(_01481_),
    .B(_01500_),
    .C(_01501_),
    .Y(_01503_));
 sky130_fd_sc_hd__a21oi_1 _08031_ (.A1(_01500_),
    .A2(_01501_),
    .B1(_01481_),
    .Y(_01504_));
 sky130_fd_sc_hd__a211oi_1 _08032_ (.A1(_01343_),
    .A2(_01347_),
    .B1(_01502_),
    .C1(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__a211o_1 _08033_ (.A1(_01343_),
    .A2(_01347_),
    .B1(_01502_),
    .C1(_01504_),
    .X(_01506_));
 sky130_fd_sc_hd__o211ai_2 _08034_ (.A1(_01502_),
    .A2(_01504_),
    .B1(_01343_),
    .C1(_01347_),
    .Y(_01507_));
 sky130_fd_sc_hd__and4_1 _08035_ (.A(_01468_),
    .B(_01469_),
    .C(_01506_),
    .D(_01507_),
    .X(_01509_));
 sky130_fd_sc_hd__a22oi_2 _08036_ (.A1(_01468_),
    .A2(_01469_),
    .B1(_01506_),
    .B2(_01507_),
    .Y(_01510_));
 sky130_fd_sc_hd__a211o_1 _08037_ (.A1(_01349_),
    .A2(_01351_),
    .B1(_01509_),
    .C1(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__o211ai_1 _08038_ (.A1(_01509_),
    .A2(_01510_),
    .B1(_01349_),
    .C1(_01351_),
    .Y(_01512_));
 sky130_fd_sc_hd__or4bb_2 _08039_ (.A(_01447_),
    .B(_01448_),
    .C_N(_01511_),
    .D_N(_01512_),
    .X(_01513_));
 sky130_fd_sc_hd__a2bb2o_1 _08040_ (.A1_N(_01447_),
    .A2_N(_01448_),
    .B1(_01511_),
    .B2(_01512_),
    .X(_01514_));
 sky130_fd_sc_hd__o211ai_2 _08041_ (.A1(_01353_),
    .A2(_01356_),
    .B1(_01513_),
    .C1(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__a211o_1 _08042_ (.A1(_01513_),
    .A2(_01514_),
    .B1(_01353_),
    .C1(_01356_),
    .X(_01516_));
 sky130_fd_sc_hd__or4bb_2 _08043_ (.A(_01407_),
    .B(_01408_),
    .C_N(_01515_),
    .D_N(_01516_),
    .X(_01517_));
 sky130_fd_sc_hd__a2bb2o_1 _08044_ (.A1_N(_01407_),
    .A2_N(_01408_),
    .B1(_01515_),
    .B2(_01516_),
    .X(_01518_));
 sky130_fd_sc_hd__o211a_1 _08045_ (.A1(_01358_),
    .A2(_01361_),
    .B1(_01517_),
    .C1(_01518_),
    .X(_01520_));
 sky130_fd_sc_hd__a211oi_1 _08046_ (.A1(_01517_),
    .A2(_01518_),
    .B1(_01358_),
    .C1(_01361_),
    .Y(_01521_));
 sky130_fd_sc_hd__a211oi_2 _08047_ (.A1(_01250_),
    .A2(_01252_),
    .B1(_01520_),
    .C1(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hd__o211a_1 _08048_ (.A1(_01520_),
    .A2(_01521_),
    .B1(_01250_),
    .C1(_01252_),
    .X(_01523_));
 sky130_fd_sc_hd__a211o_1 _08049_ (.A1(_01364_),
    .A2(_01367_),
    .B1(_01522_),
    .C1(_01523_),
    .X(_01524_));
 sky130_fd_sc_hd__o211ai_1 _08050_ (.A1(_01522_),
    .A2(_01523_),
    .B1(_01364_),
    .C1(_01367_),
    .Y(_01525_));
 sky130_fd_sc_hd__a21oi_1 _08051_ (.A1(_01524_),
    .A2(_01525_),
    .B1(_01369_),
    .Y(_01526_));
 sky130_fd_sc_hd__and3_1 _08052_ (.A(_01369_),
    .B(_01524_),
    .C(_01525_),
    .X(_01527_));
 sky130_fd_sc_hd__or2_1 _08053_ (.A(_01526_),
    .B(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__o21bai_1 _08054_ (.A1(_01221_),
    .A2(_01373_),
    .B1_N(_01372_),
    .Y(_01529_));
 sky130_fd_sc_hd__xnor2_1 _08055_ (.A(_01528_),
    .B(_01529_),
    .Y(net86));
 sky130_fd_sc_hd__nand2b_1 _08056_ (.A_N(_01401_),
    .B(_01403_),
    .Y(_01531_));
 sky130_fd_sc_hd__nand2_1 _08057_ (.A(net26),
    .B(net53),
    .Y(_01532_));
 sky130_fd_sc_hd__and4_1 _08058_ (.A(net26),
    .B(net23),
    .C(net52),
    .D(net53),
    .X(_01533_));
 sky130_fd_sc_hd__a22oi_1 _08059_ (.A1(net26),
    .A2(net52),
    .B1(net53),
    .B2(net23),
    .Y(_01534_));
 sky130_fd_sc_hd__nor2_1 _08060_ (.A(_01533_),
    .B(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__nand2_1 _08061_ (.A(net12),
    .B(net54),
    .Y(_01536_));
 sky130_fd_sc_hd__xnor2_1 _08062_ (.A(_01535_),
    .B(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__o21ba_1 _08063_ (.A1(_01377_),
    .A2(_01379_),
    .B1_N(_01375_),
    .X(_01538_));
 sky130_fd_sc_hd__nand2b_1 _08064_ (.A_N(_01538_),
    .B(_01537_),
    .Y(_01539_));
 sky130_fd_sc_hd__xnor2_1 _08065_ (.A(_01537_),
    .B(_01538_),
    .Y(_01541_));
 sky130_fd_sc_hd__nand3_1 _08066_ (.A(net1),
    .B(net56),
    .C(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__a21o_1 _08067_ (.A1(net1),
    .A2(net56),
    .B1(_01541_),
    .X(_01543_));
 sky130_fd_sc_hd__nand2_1 _08068_ (.A(_01542_),
    .B(_01543_),
    .Y(_01544_));
 sky130_fd_sc_hd__or2_1 _08069_ (.A(_01381_),
    .B(_01544_),
    .X(_01545_));
 sky130_fd_sc_hd__nand2_1 _08070_ (.A(_01381_),
    .B(_01544_),
    .Y(_01546_));
 sky130_fd_sc_hd__nand2_1 _08071_ (.A(_01545_),
    .B(_01546_),
    .Y(_01547_));
 sky130_fd_sc_hd__nor2_1 _08072_ (.A(_01386_),
    .B(_01390_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_1 _08073_ (.A(_01411_),
    .B(_01414_),
    .Y(_01549_));
 sky130_fd_sc_hd__and4_1 _08074_ (.A(net28),
    .B(net29),
    .C(net49),
    .D(net50),
    .X(_01550_));
 sky130_fd_sc_hd__a22o_1 _08075_ (.A1(net29),
    .A2(net49),
    .B1(net50),
    .B2(net28),
    .X(_01552_));
 sky130_fd_sc_hd__and2b_1 _08076_ (.A_N(_01550_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__nand2_1 _08077_ (.A(net27),
    .B(net51),
    .Y(_01554_));
 sky130_fd_sc_hd__xnor2_1 _08078_ (.A(_01553_),
    .B(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2b_1 _08079_ (.A_N(_01549_),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__xnor2_1 _08080_ (.A(_01549_),
    .B(_01555_),
    .Y(_01557_));
 sky130_fd_sc_hd__nand2b_1 _08081_ (.A_N(_01548_),
    .B(_01557_),
    .Y(_01558_));
 sky130_fd_sc_hd__xnor2_1 _08082_ (.A(_01548_),
    .B(_01557_),
    .Y(_01559_));
 sky130_fd_sc_hd__o21a_2 _08083_ (.A1(_01423_),
    .A2(_01425_),
    .B1(_01559_),
    .X(_01560_));
 sky130_fd_sc_hd__nor3_1 _08084_ (.A(_01423_),
    .B(_01425_),
    .C(_01559_),
    .Y(_01561_));
 sky130_fd_sc_hd__a211oi_4 _08085_ (.A1(_01392_),
    .A2(_01394_),
    .B1(_01560_),
    .C1(_01561_),
    .Y(_01563_));
 sky130_fd_sc_hd__o211a_1 _08086_ (.A1(_01560_),
    .A2(_01561_),
    .B1(_01392_),
    .C1(_01394_),
    .X(_01564_));
 sky130_fd_sc_hd__a211oi_2 _08087_ (.A1(_01396_),
    .A2(_01399_),
    .B1(_01563_),
    .C1(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__inv_2 _08088_ (.A(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__o211a_1 _08089_ (.A1(_01563_),
    .A2(_01564_),
    .B1(_01396_),
    .C1(_01399_),
    .X(_01567_));
 sky130_fd_sc_hd__or3_2 _08090_ (.A(_01547_),
    .B(_01565_),
    .C(_01567_),
    .X(_01568_));
 sky130_fd_sc_hd__o21ai_2 _08091_ (.A1(_01565_),
    .A2(_01567_),
    .B1(_01547_),
    .Y(_01569_));
 sky130_fd_sc_hd__o211ai_4 _08092_ (.A1(_01445_),
    .A2(_01447_),
    .B1(_01568_),
    .C1(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__a211o_1 _08093_ (.A1(_01568_),
    .A2(_01569_),
    .B1(_01445_),
    .C1(_01447_),
    .X(_01571_));
 sky130_fd_sc_hd__nand3_2 _08094_ (.A(_01531_),
    .B(_01570_),
    .C(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__a21o_1 _08095_ (.A1(_01570_),
    .A2(_01571_),
    .B1(_01531_),
    .X(_01574_));
 sky130_fd_sc_hd__nand2_1 _08096_ (.A(net32),
    .B(net47),
    .Y(_01575_));
 sky130_fd_sc_hd__and4_1 _08097_ (.A(net31),
    .B(net32),
    .C(net46),
    .D(net47),
    .X(_01576_));
 sky130_fd_sc_hd__a22o_1 _08098_ (.A1(net32),
    .A2(net46),
    .B1(net47),
    .B2(net31),
    .X(_01577_));
 sky130_fd_sc_hd__and2b_1 _08099_ (.A_N(_01576_),
    .B(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__nand2_1 _08100_ (.A(net30),
    .B(net48),
    .Y(_01579_));
 sky130_fd_sc_hd__xnor2_1 _08101_ (.A(_01578_),
    .B(_01579_),
    .Y(_01580_));
 sky130_fd_sc_hd__nand2_1 _08102_ (.A(net2),
    .B(net45),
    .Y(_01581_));
 sky130_fd_sc_hd__nand2_1 _08103_ (.A(net4),
    .B(net43),
    .Y(_01582_));
 sky130_fd_sc_hd__and4_1 _08104_ (.A(net3),
    .B(net4),
    .C(net42),
    .D(net43),
    .X(_01583_));
 sky130_fd_sc_hd__a22oi_2 _08105_ (.A1(net4),
    .A2(net42),
    .B1(net43),
    .B2(net3),
    .Y(_01585_));
 sky130_fd_sc_hd__or3_1 _08106_ (.A(_01581_),
    .B(_01583_),
    .C(_01585_),
    .X(_01586_));
 sky130_fd_sc_hd__o21ai_1 _08107_ (.A1(_01583_),
    .A2(_01585_),
    .B1(_01581_),
    .Y(_01587_));
 sky130_fd_sc_hd__o21bai_1 _08108_ (.A1(_01416_),
    .A2(_01418_),
    .B1_N(_01417_),
    .Y(_01588_));
 sky130_fd_sc_hd__and3_1 _08109_ (.A(_01586_),
    .B(_01587_),
    .C(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__a21o_1 _08110_ (.A1(_01586_),
    .A2(_01587_),
    .B1(_01588_),
    .X(_01590_));
 sky130_fd_sc_hd__and2b_1 _08111_ (.A_N(_01589_),
    .B(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__xnor2_1 _08112_ (.A(_01580_),
    .B(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__a31o_1 _08113_ (.A1(net4),
    .A2(net41),
    .A3(_01433_),
    .B1(_01430_),
    .X(_01593_));
 sky130_fd_sc_hd__o21bai_1 _08114_ (.A1(_01449_),
    .A2(_01451_),
    .B1_N(_01450_),
    .Y(_01594_));
 sky130_fd_sc_hd__nand4_1 _08115_ (.A(net6),
    .B(net7),
    .C(net39),
    .D(net40),
    .Y(_01596_));
 sky130_fd_sc_hd__a22o_1 _08116_ (.A1(net7),
    .A2(net39),
    .B1(net40),
    .B2(net6),
    .X(_01597_));
 sky130_fd_sc_hd__a22o_1 _08117_ (.A1(net5),
    .A2(net41),
    .B1(_01596_),
    .B2(_01597_),
    .X(_01598_));
 sky130_fd_sc_hd__nand4_1 _08118_ (.A(net5),
    .B(net41),
    .C(_01596_),
    .D(_01597_),
    .Y(_01599_));
 sky130_fd_sc_hd__and3_1 _08119_ (.A(_01594_),
    .B(_01598_),
    .C(_01599_),
    .X(_01600_));
 sky130_fd_sc_hd__a21o_1 _08120_ (.A1(_01598_),
    .A2(_01599_),
    .B1(_01594_),
    .X(_01601_));
 sky130_fd_sc_hd__and2b_1 _08121_ (.A_N(_01600_),
    .B(_01601_),
    .X(_01602_));
 sky130_fd_sc_hd__xnor2_1 _08122_ (.A(_01593_),
    .B(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__a21oi_1 _08123_ (.A1(_01436_),
    .A2(_01438_),
    .B1(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__and3_1 _08124_ (.A(_01436_),
    .B(_01438_),
    .C(_01603_),
    .X(_01605_));
 sky130_fd_sc_hd__nor3_1 _08125_ (.A(_01592_),
    .B(_01604_),
    .C(_01605_),
    .Y(_01607_));
 sky130_fd_sc_hd__o21a_1 _08126_ (.A1(_01604_),
    .A2(_01605_),
    .B1(_01592_),
    .X(_01608_));
 sky130_fd_sc_hd__a211oi_2 _08127_ (.A1(_01466_),
    .A2(_01468_),
    .B1(_01607_),
    .C1(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__o211a_1 _08128_ (.A1(_01607_),
    .A2(_01608_),
    .B1(_01466_),
    .C1(_01468_),
    .X(_01610_));
 sky130_fd_sc_hd__a211oi_2 _08129_ (.A1(_01440_),
    .A2(_01443_),
    .B1(_01609_),
    .C1(_01610_),
    .Y(_01611_));
 sky130_fd_sc_hd__o211a_1 _08130_ (.A1(_01609_),
    .A2(_01610_),
    .B1(_01440_),
    .C1(_01443_),
    .X(_01612_));
 sky130_fd_sc_hd__a21o_1 _08131_ (.A1(_01470_),
    .A2(_01479_),
    .B1(_01478_),
    .X(_01613_));
 sky130_fd_sc_hd__nand2_1 _08132_ (.A(net38),
    .B(net8),
    .Y(_01614_));
 sky130_fd_sc_hd__nand2_1 _08133_ (.A(net37),
    .B(net10),
    .Y(_01615_));
 sky130_fd_sc_hd__and4_1 _08134_ (.A(net36),
    .B(net37),
    .C(net9),
    .D(net10),
    .X(_01616_));
 sky130_fd_sc_hd__a22o_1 _08135_ (.A1(net37),
    .A2(net9),
    .B1(net10),
    .B2(net36),
    .X(_01618_));
 sky130_fd_sc_hd__and2b_1 _08136_ (.A_N(_01616_),
    .B(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__xnor2_1 _08137_ (.A(_01614_),
    .B(_01619_),
    .Y(_01620_));
 sky130_fd_sc_hd__nand2_1 _08138_ (.A(net35),
    .B(net11),
    .Y(_01621_));
 sky130_fd_sc_hd__nand2_1 _08139_ (.A(net34),
    .B(net14),
    .Y(_01622_));
 sky130_fd_sc_hd__and4_1 _08140_ (.A(net64),
    .B(net34),
    .C(net13),
    .D(net14),
    .X(_01623_));
 sky130_fd_sc_hd__a22oi_2 _08141_ (.A1(net34),
    .A2(net13),
    .B1(net14),
    .B2(net64),
    .Y(_01624_));
 sky130_fd_sc_hd__or3_1 _08142_ (.A(_01621_),
    .B(_01623_),
    .C(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__o21ai_1 _08143_ (.A1(_01623_),
    .A2(_01624_),
    .B1(_01621_),
    .Y(_01626_));
 sky130_fd_sc_hd__a31o_1 _08144_ (.A1(net35),
    .A2(net10),
    .A3(_01457_),
    .B1(_01456_),
    .X(_01627_));
 sky130_fd_sc_hd__nand3_2 _08145_ (.A(_01625_),
    .B(_01626_),
    .C(_01627_),
    .Y(_01629_));
 sky130_fd_sc_hd__a21o_1 _08146_ (.A1(_01625_),
    .A2(_01626_),
    .B1(_01627_),
    .X(_01630_));
 sky130_fd_sc_hd__nand3_2 _08147_ (.A(_01620_),
    .B(_01629_),
    .C(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__a21o_1 _08148_ (.A1(_01629_),
    .A2(_01630_),
    .B1(_01620_),
    .X(_01632_));
 sky130_fd_sc_hd__nand3_2 _08149_ (.A(_01613_),
    .B(_01631_),
    .C(_01632_),
    .Y(_01633_));
 sky130_fd_sc_hd__a21o_1 _08150_ (.A1(_01631_),
    .A2(_01632_),
    .B1(_01613_),
    .X(_01634_));
 sky130_fd_sc_hd__o211ai_2 _08151_ (.A1(_01461_),
    .A2(_01463_),
    .B1(_01633_),
    .C1(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__a211o_1 _08152_ (.A1(_01633_),
    .A2(_01634_),
    .B1(_01461_),
    .C1(_01463_),
    .X(_01636_));
 sky130_fd_sc_hd__nand2_1 _08153_ (.A(_01635_),
    .B(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__nand2_1 _08154_ (.A(_01473_),
    .B(_01476_),
    .Y(_01638_));
 sky130_fd_sc_hd__o21bai_1 _08155_ (.A1(_01482_),
    .A2(_01484_),
    .B1_N(_01483_),
    .Y(_01640_));
 sky130_fd_sc_hd__nand2_1 _08156_ (.A(net63),
    .B(net15),
    .Y(_01641_));
 sky130_fd_sc_hd__nand4_1 _08157_ (.A(net61),
    .B(net62),
    .C(net16),
    .D(net17),
    .Y(_01642_));
 sky130_fd_sc_hd__a22o_1 _08158_ (.A1(net62),
    .A2(net16),
    .B1(net17),
    .B2(net61),
    .X(_01643_));
 sky130_fd_sc_hd__nand3b_1 _08159_ (.A_N(_01641_),
    .B(_01642_),
    .C(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__a21bo_1 _08160_ (.A1(_01642_),
    .A2(_01643_),
    .B1_N(_01641_),
    .X(_01645_));
 sky130_fd_sc_hd__and3_1 _08161_ (.A(_01640_),
    .B(_01644_),
    .C(_01645_),
    .X(_01646_));
 sky130_fd_sc_hd__a21o_1 _08162_ (.A1(_01644_),
    .A2(_01645_),
    .B1(_01640_),
    .X(_01647_));
 sky130_fd_sc_hd__and2b_1 _08163_ (.A_N(_01646_),
    .B(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__xor2_1 _08164_ (.A(_01638_),
    .B(_01648_),
    .X(_01649_));
 sky130_fd_sc_hd__nand2_1 _08165_ (.A(net60),
    .B(net18),
    .Y(_01651_));
 sky130_fd_sc_hd__and2_1 _08166_ (.A(net59),
    .B(net20),
    .X(_01652_));
 sky130_fd_sc_hd__and4_1 _08167_ (.A(net58),
    .B(net59),
    .C(net19),
    .D(net20),
    .X(_01653_));
 sky130_fd_sc_hd__a22o_1 _08168_ (.A1(net59),
    .A2(net19),
    .B1(net20),
    .B2(net58),
    .X(_01654_));
 sky130_fd_sc_hd__and2b_1 _08169_ (.A_N(_01653_),
    .B(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__xnor2_1 _08170_ (.A(_01651_),
    .B(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__nand2_1 _08171_ (.A(net55),
    .B(net21),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_1 _08172_ (.A(net44),
    .B(net24),
    .Y(_01658_));
 sky130_fd_sc_hd__and4_1 _08173_ (.A(net33),
    .B(net44),
    .C(net22),
    .D(net24),
    .X(_01659_));
 sky130_fd_sc_hd__a22oi_2 _08174_ (.A1(net44),
    .A2(net22),
    .B1(net24),
    .B2(net33),
    .Y(_01660_));
 sky130_fd_sc_hd__nor3_1 _08175_ (.A(_01657_),
    .B(_01659_),
    .C(_01660_),
    .Y(_01662_));
 sky130_fd_sc_hd__or3_1 _08176_ (.A(_01657_),
    .B(_01659_),
    .C(_01660_),
    .X(_01663_));
 sky130_fd_sc_hd__o21ai_1 _08177_ (.A1(_01659_),
    .A2(_01660_),
    .B1(_01657_),
    .Y(_01664_));
 sky130_fd_sc_hd__a21bo_1 _08178_ (.A1(_01488_),
    .A2(_01490_),
    .B1_N(_01489_),
    .X(_01665_));
 sky130_fd_sc_hd__nand3_1 _08179_ (.A(_01663_),
    .B(_01664_),
    .C(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__a21o_1 _08180_ (.A1(_01663_),
    .A2(_01664_),
    .B1(_01665_),
    .X(_01667_));
 sky130_fd_sc_hd__nand3_1 _08181_ (.A(_01656_),
    .B(_01666_),
    .C(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__a21o_1 _08182_ (.A1(_01666_),
    .A2(_01667_),
    .B1(_01656_),
    .X(_01669_));
 sky130_fd_sc_hd__a21bo_1 _08183_ (.A1(_01487_),
    .A2(_01495_),
    .B1_N(_01494_),
    .X(_01670_));
 sky130_fd_sc_hd__nand3_4 _08184_ (.A(_01668_),
    .B(_01669_),
    .C(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__a21o_1 _08185_ (.A1(_01668_),
    .A2(_01669_),
    .B1(_01670_),
    .X(_01673_));
 sky130_fd_sc_hd__and3_1 _08186_ (.A(_01649_),
    .B(_01671_),
    .C(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__nand3_2 _08187_ (.A(_01649_),
    .B(_01671_),
    .C(_01673_),
    .Y(_01675_));
 sky130_fd_sc_hd__a21oi_1 _08188_ (.A1(_01671_),
    .A2(_01673_),
    .B1(_01649_),
    .Y(_01676_));
 sky130_fd_sc_hd__a211o_1 _08189_ (.A1(_01500_),
    .A2(_01503_),
    .B1(_01674_),
    .C1(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__o211ai_2 _08190_ (.A1(_01674_),
    .A2(_01676_),
    .B1(_01500_),
    .C1(_01503_),
    .Y(_01678_));
 sky130_fd_sc_hd__nand3b_2 _08191_ (.A_N(_01637_),
    .B(_01677_),
    .C(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hd__a21bo_1 _08192_ (.A1(_01677_),
    .A2(_01678_),
    .B1_N(_01637_),
    .X(_01680_));
 sky130_fd_sc_hd__o211a_1 _08193_ (.A1(_01505_),
    .A2(_01509_),
    .B1(_01679_),
    .C1(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__a211oi_2 _08194_ (.A1(_01679_),
    .A2(_01680_),
    .B1(_01505_),
    .C1(_01509_),
    .Y(_01682_));
 sky130_fd_sc_hd__nor4_2 _08195_ (.A(_01611_),
    .B(_01612_),
    .C(_01681_),
    .D(_01682_),
    .Y(_01684_));
 sky130_fd_sc_hd__o22a_1 _08196_ (.A1(_01611_),
    .A2(_01612_),
    .B1(_01681_),
    .B2(_01682_),
    .X(_01685_));
 sky130_fd_sc_hd__a211oi_1 _08197_ (.A1(_01511_),
    .A2(_01513_),
    .B1(_01684_),
    .C1(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__a211o_1 _08198_ (.A1(_01511_),
    .A2(_01513_),
    .B1(_01684_),
    .C1(_01685_),
    .X(_01687_));
 sky130_fd_sc_hd__o211ai_1 _08199_ (.A1(_01684_),
    .A2(_01685_),
    .B1(_01511_),
    .C1(_01513_),
    .Y(_01688_));
 sky130_fd_sc_hd__and4_1 _08200_ (.A(_01572_),
    .B(_01574_),
    .C(_01687_),
    .D(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__a22oi_2 _08201_ (.A1(_01572_),
    .A2(_01574_),
    .B1(_01687_),
    .B2(_01688_),
    .Y(_01690_));
 sky130_fd_sc_hd__a211o_1 _08202_ (.A1(_01515_),
    .A2(_01517_),
    .B1(_01689_),
    .C1(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__o211ai_2 _08203_ (.A1(_01689_),
    .A2(_01690_),
    .B1(_01515_),
    .C1(_01517_),
    .Y(_01692_));
 sky130_fd_sc_hd__o211ai_2 _08204_ (.A1(_01405_),
    .A2(_01407_),
    .B1(_01691_),
    .C1(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__a211o_1 _08205_ (.A1(_01691_),
    .A2(_01692_),
    .B1(_01405_),
    .C1(_01407_),
    .X(_01694_));
 sky130_fd_sc_hd__o211a_1 _08206_ (.A1(_01520_),
    .A2(_01522_),
    .B1(_01693_),
    .C1(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__a211oi_1 _08207_ (.A1(_01693_),
    .A2(_01694_),
    .B1(_01520_),
    .C1(_01522_),
    .Y(_01696_));
 sky130_fd_sc_hd__nor2_1 _08208_ (.A(_01695_),
    .B(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__and2b_1 _08209_ (.A_N(_01524_),
    .B(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__xnor2_1 _08210_ (.A(_01524_),
    .B(_01697_),
    .Y(_01699_));
 sky130_fd_sc_hd__nor2_1 _08211_ (.A(_01372_),
    .B(_01527_),
    .Y(_01700_));
 sky130_fd_sc_hd__nor2_1 _08212_ (.A(_01526_),
    .B(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__or4_1 _08213_ (.A(_01372_),
    .B(_01373_),
    .C(_01526_),
    .D(_01527_),
    .X(_01702_));
 sky130_fd_sc_hd__o21ba_1 _08214_ (.A1(_01221_),
    .A2(_01702_),
    .B1_N(_01701_),
    .X(_01703_));
 sky130_fd_sc_hd__and2b_1 _08215_ (.A_N(_01703_),
    .B(_01699_),
    .X(_01705_));
 sky130_fd_sc_hd__xnor2_1 _08216_ (.A(_01699_),
    .B(_01703_),
    .Y(net88));
 sky130_fd_sc_hd__and4_1 _08217_ (.A(net28),
    .B(net27),
    .C(net51),
    .D(net52),
    .X(_01706_));
 sky130_fd_sc_hd__a22o_1 _08218_ (.A1(net28),
    .A2(net51),
    .B1(net52),
    .B2(net27),
    .X(_01707_));
 sky130_fd_sc_hd__and2b_1 _08219_ (.A_N(_01706_),
    .B(_01707_),
    .X(_01708_));
 sky130_fd_sc_hd__xnor2_1 _08220_ (.A(_01532_),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__o21ba_1 _08221_ (.A1(_01534_),
    .A2(_01536_),
    .B1_N(_01533_),
    .X(_01710_));
 sky130_fd_sc_hd__and2b_1 _08222_ (.A_N(_01710_),
    .B(_01709_),
    .X(_01711_));
 sky130_fd_sc_hd__xnor2_1 _08223_ (.A(_01709_),
    .B(_01710_),
    .Y(_01712_));
 sky130_fd_sc_hd__nand2_1 _08224_ (.A(net23),
    .B(net56),
    .Y(_01713_));
 sky130_fd_sc_hd__nor2_1 _08225_ (.A(_01536_),
    .B(_01713_),
    .Y(_01715_));
 sky130_fd_sc_hd__or2_1 _08226_ (.A(_01536_),
    .B(_01713_),
    .X(_01716_));
 sky130_fd_sc_hd__a22o_1 _08227_ (.A1(net23),
    .A2(net54),
    .B1(net56),
    .B2(net12),
    .X(_01717_));
 sky130_fd_sc_hd__o2bb2a_1 _08228_ (.A1_N(_01716_),
    .A2_N(_01717_),
    .B1(net1),
    .B2(_00287_),
    .X(_01718_));
 sky130_fd_sc_hd__and4b_1 _08229_ (.A_N(net1),
    .B(net57),
    .C(_01716_),
    .D(_01717_),
    .X(_01719_));
 sky130_fd_sc_hd__nor2_1 _08230_ (.A(_01718_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__nor2_1 _08231_ (.A(_01712_),
    .B(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__and2_1 _08232_ (.A(_01712_),
    .B(_01720_),
    .X(_01722_));
 sky130_fd_sc_hd__or2_1 _08233_ (.A(_01721_),
    .B(_01722_),
    .X(_01723_));
 sky130_fd_sc_hd__a21o_1 _08234_ (.A1(_01539_),
    .A2(_01542_),
    .B1(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__nand3_1 _08235_ (.A(_01539_),
    .B(_01542_),
    .C(_01723_),
    .Y(_01726_));
 sky130_fd_sc_hd__a21o_1 _08236_ (.A1(_01580_),
    .A2(_01590_),
    .B1(_01589_),
    .X(_01727_));
 sky130_fd_sc_hd__a31o_1 _08237_ (.A1(net27),
    .A2(net51),
    .A3(_01552_),
    .B1(_01550_),
    .X(_01728_));
 sky130_fd_sc_hd__a31o_1 _08238_ (.A1(net30),
    .A2(net48),
    .A3(_01577_),
    .B1(_01576_),
    .X(_01729_));
 sky130_fd_sc_hd__nand4_1 _08239_ (.A(net30),
    .B(net31),
    .C(net48),
    .D(net49),
    .Y(_01730_));
 sky130_fd_sc_hd__a22o_1 _08240_ (.A1(net31),
    .A2(net48),
    .B1(net49),
    .B2(net30),
    .X(_01731_));
 sky130_fd_sc_hd__a22o_1 _08241_ (.A1(net29),
    .A2(net50),
    .B1(_01730_),
    .B2(_01731_),
    .X(_01732_));
 sky130_fd_sc_hd__nand4_1 _08242_ (.A(net29),
    .B(net50),
    .C(_01730_),
    .D(_01731_),
    .Y(_01733_));
 sky130_fd_sc_hd__nand3_1 _08243_ (.A(_01729_),
    .B(_01732_),
    .C(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__a21o_1 _08244_ (.A1(_01732_),
    .A2(_01733_),
    .B1(_01729_),
    .X(_01735_));
 sky130_fd_sc_hd__nand3_1 _08245_ (.A(_01728_),
    .B(_01734_),
    .C(_01735_),
    .Y(_01737_));
 sky130_fd_sc_hd__a21o_1 _08246_ (.A1(_01734_),
    .A2(_01735_),
    .B1(_01728_),
    .X(_01738_));
 sky130_fd_sc_hd__and3_1 _08247_ (.A(_01727_),
    .B(_01737_),
    .C(_01738_),
    .X(_01739_));
 sky130_fd_sc_hd__a21oi_2 _08248_ (.A1(_01737_),
    .A2(_01738_),
    .B1(_01727_),
    .Y(_01740_));
 sky130_fd_sc_hd__a211oi_2 _08249_ (.A1(_01556_),
    .A2(_01558_),
    .B1(_01739_),
    .C1(_01740_),
    .Y(_01741_));
 sky130_fd_sc_hd__inv_2 _08250_ (.A(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__o211ai_2 _08251_ (.A1(_01739_),
    .A2(_01740_),
    .B1(_01556_),
    .C1(_01558_),
    .Y(_01743_));
 sky130_fd_sc_hd__o211ai_2 _08252_ (.A1(_01560_),
    .A2(_01563_),
    .B1(_01742_),
    .C1(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__a211o_1 _08253_ (.A1(_01742_),
    .A2(_01743_),
    .B1(_01560_),
    .C1(_01563_),
    .X(_01745_));
 sky130_fd_sc_hd__nand4_1 _08254_ (.A(_01724_),
    .B(_01726_),
    .C(_01744_),
    .D(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__a22o_1 _08255_ (.A1(_01724_),
    .A2(_01726_),
    .B1(_01744_),
    .B2(_01745_),
    .X(_01748_));
 sky130_fd_sc_hd__o211a_1 _08256_ (.A1(_01609_),
    .A2(_01611_),
    .B1(_01746_),
    .C1(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__a211oi_1 _08257_ (.A1(_01746_),
    .A2(_01748_),
    .B1(_01609_),
    .C1(_01611_),
    .Y(_01750_));
 sky130_fd_sc_hd__a211oi_1 _08258_ (.A1(_01566_),
    .A2(_01568_),
    .B1(_01749_),
    .C1(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__o211a_1 _08259_ (.A1(_01749_),
    .A2(_01750_),
    .B1(_01566_),
    .C1(_01568_),
    .X(_01752_));
 sky130_fd_sc_hd__nand2_1 _08260_ (.A(_01633_),
    .B(_01635_),
    .Y(_01753_));
 sky130_fd_sc_hd__and4_1 _08261_ (.A(net2),
    .B(net3),
    .C(net45),
    .D(net46),
    .X(_01754_));
 sky130_fd_sc_hd__a22o_1 _08262_ (.A1(net3),
    .A2(net45),
    .B1(net46),
    .B2(net2),
    .X(_01755_));
 sky130_fd_sc_hd__and2b_1 _08263_ (.A_N(_01754_),
    .B(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__xnor2_1 _08264_ (.A(_01575_),
    .B(_01756_),
    .Y(_01757_));
 sky130_fd_sc_hd__and4_1 _08265_ (.A(net5),
    .B(net6),
    .C(net41),
    .D(net42),
    .X(_01759_));
 sky130_fd_sc_hd__a22oi_2 _08266_ (.A1(net6),
    .A2(net41),
    .B1(net42),
    .B2(net5),
    .Y(_01760_));
 sky130_fd_sc_hd__or3_1 _08267_ (.A(_01582_),
    .B(_01759_),
    .C(_01760_),
    .X(_01761_));
 sky130_fd_sc_hd__o21ai_1 _08268_ (.A1(_01759_),
    .A2(_01760_),
    .B1(_01582_),
    .Y(_01762_));
 sky130_fd_sc_hd__o21bai_1 _08269_ (.A1(_01581_),
    .A2(_01585_),
    .B1_N(_01583_),
    .Y(_01763_));
 sky130_fd_sc_hd__and3_1 _08270_ (.A(_01761_),
    .B(_01762_),
    .C(_01763_),
    .X(_01764_));
 sky130_fd_sc_hd__a21o_1 _08271_ (.A1(_01761_),
    .A2(_01762_),
    .B1(_01763_),
    .X(_01765_));
 sky130_fd_sc_hd__and2b_1 _08272_ (.A_N(_01764_),
    .B(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__xnor2_1 _08273_ (.A(_01757_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__nand2_1 _08274_ (.A(_01596_),
    .B(_01599_),
    .Y(_01768_));
 sky130_fd_sc_hd__a31o_1 _08275_ (.A1(net38),
    .A2(net8),
    .A3(_01618_),
    .B1(_01616_),
    .X(_01770_));
 sky130_fd_sc_hd__nand4_1 _08276_ (.A(net38),
    .B(net39),
    .C(net8),
    .D(net9),
    .Y(_01771_));
 sky130_fd_sc_hd__a22o_1 _08277_ (.A1(net39),
    .A2(net8),
    .B1(net9),
    .B2(net38),
    .X(_01772_));
 sky130_fd_sc_hd__a22o_1 _08278_ (.A1(net7),
    .A2(net40),
    .B1(_01771_),
    .B2(_01772_),
    .X(_01773_));
 sky130_fd_sc_hd__nand4_1 _08279_ (.A(net7),
    .B(net40),
    .C(_01771_),
    .D(_01772_),
    .Y(_01774_));
 sky130_fd_sc_hd__nand3_1 _08280_ (.A(_01770_),
    .B(_01773_),
    .C(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__a21o_1 _08281_ (.A1(_01773_),
    .A2(_01774_),
    .B1(_01770_),
    .X(_01776_));
 sky130_fd_sc_hd__nand3_1 _08282_ (.A(_01768_),
    .B(_01775_),
    .C(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__a21o_1 _08283_ (.A1(_01775_),
    .A2(_01776_),
    .B1(_01768_),
    .X(_01778_));
 sky130_fd_sc_hd__a21o_1 _08284_ (.A1(_01593_),
    .A2(_01601_),
    .B1(_01600_),
    .X(_01779_));
 sky130_fd_sc_hd__and3_1 _08285_ (.A(_01777_),
    .B(_01778_),
    .C(_01779_),
    .X(_01781_));
 sky130_fd_sc_hd__a21oi_1 _08286_ (.A1(_01777_),
    .A2(_01778_),
    .B1(_01779_),
    .Y(_01782_));
 sky130_fd_sc_hd__nor3_1 _08287_ (.A(_01767_),
    .B(_01781_),
    .C(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__o21a_1 _08288_ (.A1(_01781_),
    .A2(_01782_),
    .B1(_01767_),
    .X(_01784_));
 sky130_fd_sc_hd__nor2_1 _08289_ (.A(_01783_),
    .B(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__a211o_1 _08290_ (.A1(_01633_),
    .A2(_01635_),
    .B1(_01783_),
    .C1(_01784_),
    .X(_01786_));
 sky130_fd_sc_hd__o211ai_1 _08291_ (.A1(_01783_),
    .A2(_01784_),
    .B1(_01633_),
    .C1(_01635_),
    .Y(_01787_));
 sky130_fd_sc_hd__o211a_1 _08292_ (.A1(_01604_),
    .A2(_01607_),
    .B1(_01786_),
    .C1(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__a211oi_1 _08293_ (.A1(_01786_),
    .A2(_01787_),
    .B1(_01604_),
    .C1(_01607_),
    .Y(_01789_));
 sky130_fd_sc_hd__a21o_1 _08294_ (.A1(_01638_),
    .A2(_01647_),
    .B1(_01646_),
    .X(_01790_));
 sky130_fd_sc_hd__and4_1 _08295_ (.A(net35),
    .B(net36),
    .C(net11),
    .D(net13),
    .X(_01792_));
 sky130_fd_sc_hd__a22o_1 _08296_ (.A1(net36),
    .A2(net11),
    .B1(net13),
    .B2(net35),
    .X(_01793_));
 sky130_fd_sc_hd__and2b_1 _08297_ (.A_N(_01792_),
    .B(_01793_),
    .X(_01794_));
 sky130_fd_sc_hd__xnor2_1 _08298_ (.A(_01615_),
    .B(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__and4_1 _08299_ (.A(net63),
    .B(net64),
    .C(net15),
    .D(net16),
    .X(_01796_));
 sky130_fd_sc_hd__a22oi_2 _08300_ (.A1(net64),
    .A2(net15),
    .B1(net16),
    .B2(net63),
    .Y(_01797_));
 sky130_fd_sc_hd__or3_1 _08301_ (.A(_01622_),
    .B(_01796_),
    .C(_01797_),
    .X(_01798_));
 sky130_fd_sc_hd__o21ai_1 _08302_ (.A1(_01796_),
    .A2(_01797_),
    .B1(_01622_),
    .Y(_01799_));
 sky130_fd_sc_hd__o21bai_1 _08303_ (.A1(_01621_),
    .A2(_01624_),
    .B1_N(_01623_),
    .Y(_01800_));
 sky130_fd_sc_hd__nand3_1 _08304_ (.A(_01798_),
    .B(_01799_),
    .C(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__a21o_1 _08305_ (.A1(_01798_),
    .A2(_01799_),
    .B1(_01800_),
    .X(_01803_));
 sky130_fd_sc_hd__nand3_1 _08306_ (.A(_01795_),
    .B(_01801_),
    .C(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__a21o_1 _08307_ (.A1(_01801_),
    .A2(_01803_),
    .B1(_01795_),
    .X(_01805_));
 sky130_fd_sc_hd__and3_1 _08308_ (.A(_01790_),
    .B(_01804_),
    .C(_01805_),
    .X(_01806_));
 sky130_fd_sc_hd__nand3_1 _08309_ (.A(_01790_),
    .B(_01804_),
    .C(_01805_),
    .Y(_01807_));
 sky130_fd_sc_hd__a21oi_1 _08310_ (.A1(_01804_),
    .A2(_01805_),
    .B1(_01790_),
    .Y(_01808_));
 sky130_fd_sc_hd__a211o_1 _08311_ (.A1(_01629_),
    .A2(_01631_),
    .B1(_01806_),
    .C1(_01808_),
    .X(_01809_));
 sky130_fd_sc_hd__o211ai_1 _08312_ (.A1(_01806_),
    .A2(_01808_),
    .B1(_01629_),
    .C1(_01631_),
    .Y(_01810_));
 sky130_fd_sc_hd__nand2_1 _08313_ (.A(_01809_),
    .B(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__nand2_1 _08314_ (.A(_01642_),
    .B(_01644_),
    .Y(_01812_));
 sky130_fd_sc_hd__a31o_1 _08315_ (.A1(net60),
    .A2(net18),
    .A3(_01654_),
    .B1(_01653_),
    .X(_01814_));
 sky130_fd_sc_hd__a22o_1 _08316_ (.A1(net61),
    .A2(net18),
    .B1(net19),
    .B2(net60),
    .X(_01815_));
 sky130_fd_sc_hd__nand4_1 _08317_ (.A(net60),
    .B(net61),
    .C(net18),
    .D(net19),
    .Y(_01816_));
 sky130_fd_sc_hd__a22o_1 _08318_ (.A1(net62),
    .A2(net17),
    .B1(_01815_),
    .B2(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__nand4_1 _08319_ (.A(net62),
    .B(net17),
    .C(_01815_),
    .D(_01816_),
    .Y(_01818_));
 sky130_fd_sc_hd__and3_1 _08320_ (.A(_01814_),
    .B(_01817_),
    .C(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__a21o_1 _08321_ (.A1(_01817_),
    .A2(_01818_),
    .B1(_01814_),
    .X(_01820_));
 sky130_fd_sc_hd__and2b_1 _08322_ (.A_N(_01819_),
    .B(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__xor2_1 _08323_ (.A(_01812_),
    .B(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__and3_1 _08324_ (.A(net55),
    .B(net58),
    .C(net22),
    .X(_01823_));
 sky130_fd_sc_hd__a22o_1 _08325_ (.A1(net58),
    .A2(net21),
    .B1(net22),
    .B2(net55),
    .X(_01825_));
 sky130_fd_sc_hd__a21bo_1 _08326_ (.A1(net21),
    .A2(_01823_),
    .B1_N(_01825_),
    .X(_01826_));
 sky130_fd_sc_hd__xnor2_1 _08327_ (.A(_01652_),
    .B(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__a21oi_1 _08328_ (.A1(net33),
    .A2(net25),
    .B1(net57),
    .Y(_01828_));
 sky130_fd_sc_hd__and3_1 _08329_ (.A(net33),
    .B(net57),
    .C(net25),
    .X(_01829_));
 sky130_fd_sc_hd__or3_1 _08330_ (.A(_01658_),
    .B(_01828_),
    .C(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__o21ai_1 _08331_ (.A1(_01828_),
    .A2(_01829_),
    .B1(_01658_),
    .Y(_01831_));
 sky130_fd_sc_hd__o211ai_2 _08332_ (.A1(_01659_),
    .A2(_01662_),
    .B1(_01830_),
    .C1(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__a211o_1 _08333_ (.A1(_01830_),
    .A2(_01831_),
    .B1(_01659_),
    .C1(_01662_),
    .X(_01833_));
 sky130_fd_sc_hd__nand3_1 _08334_ (.A(_01827_),
    .B(_01832_),
    .C(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__a21o_1 _08335_ (.A1(_01832_),
    .A2(_01833_),
    .B1(_01827_),
    .X(_01836_));
 sky130_fd_sc_hd__a21bo_1 _08336_ (.A1(_01656_),
    .A2(_01667_),
    .B1_N(_01666_),
    .X(_01837_));
 sky130_fd_sc_hd__nand3_2 _08337_ (.A(_01834_),
    .B(_01836_),
    .C(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__a21o_1 _08338_ (.A1(_01834_),
    .A2(_01836_),
    .B1(_01837_),
    .X(_01839_));
 sky130_fd_sc_hd__and3_1 _08339_ (.A(_01822_),
    .B(_01838_),
    .C(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__nand3_1 _08340_ (.A(_01822_),
    .B(_01838_),
    .C(_01839_),
    .Y(_01841_));
 sky130_fd_sc_hd__a21oi_2 _08341_ (.A1(_01838_),
    .A2(_01839_),
    .B1(_01822_),
    .Y(_01842_));
 sky130_fd_sc_hd__a211oi_4 _08342_ (.A1(_01671_),
    .A2(_01675_),
    .B1(_01840_),
    .C1(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__o211a_1 _08343_ (.A1(_01840_),
    .A2(_01842_),
    .B1(_01671_),
    .C1(_01675_),
    .X(_01844_));
 sky130_fd_sc_hd__nor3_2 _08344_ (.A(_01811_),
    .B(_01843_),
    .C(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__o21a_1 _08345_ (.A1(_01843_),
    .A2(_01844_),
    .B1(_01811_),
    .X(_01847_));
 sky130_fd_sc_hd__a211o_1 _08346_ (.A1(_01677_),
    .A2(_01679_),
    .B1(_01845_),
    .C1(_01847_),
    .X(_01848_));
 sky130_fd_sc_hd__o211ai_1 _08347_ (.A1(_01845_),
    .A2(_01847_),
    .B1(_01677_),
    .C1(_01679_),
    .Y(_01849_));
 sky130_fd_sc_hd__or4bb_2 _08348_ (.A(_01788_),
    .B(_01789_),
    .C_N(_01848_),
    .D_N(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__a2bb2o_1 _08349_ (.A1_N(_01788_),
    .A2_N(_01789_),
    .B1(_01848_),
    .B2(_01849_),
    .X(_01851_));
 sky130_fd_sc_hd__o211ai_2 _08350_ (.A1(_01681_),
    .A2(_01684_),
    .B1(_01850_),
    .C1(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__a211o_1 _08351_ (.A1(_01850_),
    .A2(_01851_),
    .B1(_01681_),
    .C1(_01684_),
    .X(_01853_));
 sky130_fd_sc_hd__or4bb_2 _08352_ (.A(_01751_),
    .B(_01752_),
    .C_N(_01852_),
    .D_N(_01853_),
    .X(_01854_));
 sky130_fd_sc_hd__a2bb2o_1 _08353_ (.A1_N(_01751_),
    .A2_N(_01752_),
    .B1(_01852_),
    .B2(_01853_),
    .X(_01855_));
 sky130_fd_sc_hd__o211a_2 _08354_ (.A1(_01686_),
    .A2(_01689_),
    .B1(_01854_),
    .C1(_01855_),
    .X(_01856_));
 sky130_fd_sc_hd__a211oi_2 _08355_ (.A1(_01854_),
    .A2(_01855_),
    .B1(_01686_),
    .C1(_01689_),
    .Y(_01858_));
 sky130_fd_sc_hd__a211oi_4 _08356_ (.A1(_01570_),
    .A2(_01572_),
    .B1(_01856_),
    .C1(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__o211a_1 _08357_ (.A1(_01856_),
    .A2(_01858_),
    .B1(_01570_),
    .C1(_01572_),
    .X(_01860_));
 sky130_fd_sc_hd__a211oi_1 _08358_ (.A1(_01691_),
    .A2(_01693_),
    .B1(_01859_),
    .C1(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__o211a_1 _08359_ (.A1(_01859_),
    .A2(_01860_),
    .B1(_01691_),
    .C1(_01693_),
    .X(_01862_));
 sky130_fd_sc_hd__or3_1 _08360_ (.A(_01545_),
    .B(_01861_),
    .C(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__o21ai_1 _08361_ (.A1(_01861_),
    .A2(_01862_),
    .B1(_01545_),
    .Y(_01864_));
 sky130_fd_sc_hd__a21oi_1 _08362_ (.A1(_01863_),
    .A2(_01864_),
    .B1(_01695_),
    .Y(_01865_));
 sky130_fd_sc_hd__a21o_1 _08363_ (.A1(_01863_),
    .A2(_01864_),
    .B1(_01695_),
    .X(_01866_));
 sky130_fd_sc_hd__and3_1 _08364_ (.A(_01695_),
    .B(_01863_),
    .C(_01864_),
    .X(_01867_));
 sky130_fd_sc_hd__nor2_1 _08365_ (.A(_01865_),
    .B(_01867_),
    .Y(_01869_));
 sky130_fd_sc_hd__nor2_1 _08366_ (.A(_01698_),
    .B(_01705_),
    .Y(_01870_));
 sky130_fd_sc_hd__xnor2_1 _08367_ (.A(_01869_),
    .B(_01870_),
    .Y(net89));
 sky130_fd_sc_hd__or2_1 _08368_ (.A(_01749_),
    .B(_01751_),
    .X(_01871_));
 sky130_fd_sc_hd__nand2_1 _08369_ (.A(_01744_),
    .B(_01746_),
    .Y(_01872_));
 sky130_fd_sc_hd__a21oi_1 _08370_ (.A1(_01753_),
    .A2(_01785_),
    .B1(_01788_),
    .Y(_01873_));
 sky130_fd_sc_hd__nor3_1 _08371_ (.A(net12),
    .B(_00287_),
    .C(_01713_),
    .Y(_01874_));
 sky130_fd_sc_hd__inv_2 _08372_ (.A(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hd__o21a_1 _08373_ (.A1(net12),
    .A2(_00287_),
    .B1(_01713_),
    .X(_01876_));
 sky130_fd_sc_hd__nor2_1 _08374_ (.A(_01874_),
    .B(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__and4_1 _08375_ (.A(net28),
    .B(net27),
    .C(net52),
    .D(net53),
    .X(_01879_));
 sky130_fd_sc_hd__a22o_1 _08376_ (.A1(net28),
    .A2(net52),
    .B1(net53),
    .B2(net27),
    .X(_01880_));
 sky130_fd_sc_hd__and2b_1 _08377_ (.A_N(_01879_),
    .B(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__nand2_1 _08378_ (.A(net26),
    .B(net54),
    .Y(_01882_));
 sky130_fd_sc_hd__xnor2_1 _08379_ (.A(_01881_),
    .B(_01882_),
    .Y(_01883_));
 sky130_fd_sc_hd__a31o_1 _08380_ (.A1(net26),
    .A2(net53),
    .A3(_01707_),
    .B1(_01706_),
    .X(_01884_));
 sky130_fd_sc_hd__nand2_1 _08381_ (.A(_01883_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__xor2_1 _08382_ (.A(_01883_),
    .B(_01884_),
    .X(_01886_));
 sky130_fd_sc_hd__nand2_1 _08383_ (.A(_01877_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__xor2_1 _08384_ (.A(_01877_),
    .B(_01886_),
    .X(_01888_));
 sky130_fd_sc_hd__o21ai_1 _08385_ (.A1(_01711_),
    .A2(_01722_),
    .B1(_01888_),
    .Y(_01890_));
 sky130_fd_sc_hd__or3_1 _08386_ (.A(_01711_),
    .B(_01722_),
    .C(_01888_),
    .X(_01891_));
 sky130_fd_sc_hd__o211ai_1 _08387_ (.A1(_01715_),
    .A2(_01719_),
    .B1(_01890_),
    .C1(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__a211o_1 _08388_ (.A1(_01890_),
    .A2(_01891_),
    .B1(_01715_),
    .C1(_01719_),
    .X(_01893_));
 sky130_fd_sc_hd__nand2_1 _08389_ (.A(_01892_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__a21o_1 _08390_ (.A1(_01757_),
    .A2(_01765_),
    .B1(_01764_),
    .X(_01895_));
 sky130_fd_sc_hd__nand2_1 _08391_ (.A(_01730_),
    .B(_01733_),
    .Y(_01896_));
 sky130_fd_sc_hd__a31o_1 _08392_ (.A1(net32),
    .A2(net47),
    .A3(_01755_),
    .B1(_01754_),
    .X(_01897_));
 sky130_fd_sc_hd__nand4_1 _08393_ (.A(net30),
    .B(net31),
    .C(net49),
    .D(net50),
    .Y(_01898_));
 sky130_fd_sc_hd__a22o_1 _08394_ (.A1(net31),
    .A2(net49),
    .B1(net50),
    .B2(net30),
    .X(_01899_));
 sky130_fd_sc_hd__a22o_1 _08395_ (.A1(net29),
    .A2(net51),
    .B1(_01898_),
    .B2(_01899_),
    .X(_01901_));
 sky130_fd_sc_hd__nand4_1 _08396_ (.A(net29),
    .B(net51),
    .C(_01898_),
    .D(_01899_),
    .Y(_01902_));
 sky130_fd_sc_hd__nand3_1 _08397_ (.A(_01897_),
    .B(_01901_),
    .C(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__a21o_1 _08398_ (.A1(_01901_),
    .A2(_01902_),
    .B1(_01897_),
    .X(_01904_));
 sky130_fd_sc_hd__nand3_1 _08399_ (.A(_01896_),
    .B(_01903_),
    .C(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__a21o_1 _08400_ (.A1(_01903_),
    .A2(_01904_),
    .B1(_01896_),
    .X(_01906_));
 sky130_fd_sc_hd__and3_1 _08401_ (.A(_01895_),
    .B(_01905_),
    .C(_01906_),
    .X(_01907_));
 sky130_fd_sc_hd__a21oi_1 _08402_ (.A1(_01905_),
    .A2(_01906_),
    .B1(_01895_),
    .Y(_01908_));
 sky130_fd_sc_hd__a211o_1 _08403_ (.A1(_01734_),
    .A2(_01737_),
    .B1(_01907_),
    .C1(_01908_),
    .X(_01909_));
 sky130_fd_sc_hd__o211ai_1 _08404_ (.A1(_01907_),
    .A2(_01908_),
    .B1(_01734_),
    .C1(_01737_),
    .Y(_01910_));
 sky130_fd_sc_hd__o211a_1 _08405_ (.A1(_01739_),
    .A2(_01741_),
    .B1(_01909_),
    .C1(_01910_),
    .X(_01912_));
 sky130_fd_sc_hd__a211oi_1 _08406_ (.A1(_01909_),
    .A2(_01910_),
    .B1(_01739_),
    .C1(_01741_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _08407_ (.A(_01912_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__xor2_1 _08408_ (.A(_01894_),
    .B(_01914_),
    .X(_01915_));
 sky130_fd_sc_hd__nor2_1 _08409_ (.A(_01873_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__xor2_1 _08410_ (.A(_01873_),
    .B(_01915_),
    .X(_01917_));
 sky130_fd_sc_hd__xor2_1 _08411_ (.A(_01872_),
    .B(_01917_),
    .X(_01918_));
 sky130_fd_sc_hd__nor2_1 _08412_ (.A(_01781_),
    .B(_01783_),
    .Y(_01919_));
 sky130_fd_sc_hd__and4_1 _08413_ (.A(net2),
    .B(net3),
    .C(net46),
    .D(net47),
    .X(_01920_));
 sky130_fd_sc_hd__a22o_1 _08414_ (.A1(net3),
    .A2(net46),
    .B1(net47),
    .B2(net2),
    .X(_01921_));
 sky130_fd_sc_hd__and2b_1 _08415_ (.A_N(_01920_),
    .B(_01921_),
    .X(_01923_));
 sky130_fd_sc_hd__nand2_1 _08416_ (.A(net32),
    .B(net48),
    .Y(_01924_));
 sky130_fd_sc_hd__xnor2_1 _08417_ (.A(_01923_),
    .B(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand4_1 _08418_ (.A(net5),
    .B(net6),
    .C(net42),
    .D(net43),
    .Y(_01926_));
 sky130_fd_sc_hd__a22o_1 _08419_ (.A1(net6),
    .A2(net42),
    .B1(net43),
    .B2(net5),
    .X(_01927_));
 sky130_fd_sc_hd__and2_1 _08420_ (.A(net4),
    .B(net45),
    .X(_01928_));
 sky130_fd_sc_hd__a21o_1 _08421_ (.A1(_01926_),
    .A2(_01927_),
    .B1(_01928_),
    .X(_01929_));
 sky130_fd_sc_hd__nand3_1 _08422_ (.A(_01926_),
    .B(_01927_),
    .C(_01928_),
    .Y(_01930_));
 sky130_fd_sc_hd__o21bai_1 _08423_ (.A1(_01582_),
    .A2(_01760_),
    .B1_N(_01759_),
    .Y(_01931_));
 sky130_fd_sc_hd__and3_1 _08424_ (.A(_01929_),
    .B(_01930_),
    .C(_01931_),
    .X(_01932_));
 sky130_fd_sc_hd__a21o_1 _08425_ (.A1(_01929_),
    .A2(_01930_),
    .B1(_01931_),
    .X(_01934_));
 sky130_fd_sc_hd__and2b_1 _08426_ (.A_N(_01932_),
    .B(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__xnor2_1 _08427_ (.A(_01925_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__nand2_1 _08428_ (.A(_01771_),
    .B(_01774_),
    .Y(_01937_));
 sky130_fd_sc_hd__a31o_1 _08429_ (.A1(net37),
    .A2(net10),
    .A3(_01793_),
    .B1(_01792_),
    .X(_01938_));
 sky130_fd_sc_hd__nand4_1 _08430_ (.A(net39),
    .B(net8),
    .C(net40),
    .D(net9),
    .Y(_01939_));
 sky130_fd_sc_hd__a22o_1 _08431_ (.A1(net8),
    .A2(net40),
    .B1(net9),
    .B2(net39),
    .X(_01940_));
 sky130_fd_sc_hd__a22o_1 _08432_ (.A1(net7),
    .A2(net41),
    .B1(_01939_),
    .B2(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__nand4_1 _08433_ (.A(net7),
    .B(net41),
    .C(_01939_),
    .D(_01940_),
    .Y(_01942_));
 sky130_fd_sc_hd__nand3_1 _08434_ (.A(_01938_),
    .B(_01941_),
    .C(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__a21o_1 _08435_ (.A1(_01941_),
    .A2(_01942_),
    .B1(_01938_),
    .X(_01945_));
 sky130_fd_sc_hd__nand3_1 _08436_ (.A(_01937_),
    .B(_01943_),
    .C(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__a21o_1 _08437_ (.A1(_01943_),
    .A2(_01945_),
    .B1(_01937_),
    .X(_01947_));
 sky130_fd_sc_hd__a21bo_1 _08438_ (.A1(_01768_),
    .A2(_01776_),
    .B1_N(_01775_),
    .X(_01948_));
 sky130_fd_sc_hd__and3_1 _08439_ (.A(_01946_),
    .B(_01947_),
    .C(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__a21oi_1 _08440_ (.A1(_01946_),
    .A2(_01947_),
    .B1(_01948_),
    .Y(_01950_));
 sky130_fd_sc_hd__nor3_1 _08441_ (.A(_01936_),
    .B(_01949_),
    .C(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__o21a_1 _08442_ (.A1(_01949_),
    .A2(_01950_),
    .B1(_01936_),
    .X(_01952_));
 sky130_fd_sc_hd__a211oi_1 _08443_ (.A1(_01807_),
    .A2(_01809_),
    .B1(_01951_),
    .C1(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__o211a_1 _08444_ (.A1(_01951_),
    .A2(_01952_),
    .B1(_01807_),
    .C1(_01809_),
    .X(_01954_));
 sky130_fd_sc_hd__nor2_1 _08445_ (.A(_01953_),
    .B(_01954_),
    .Y(_01956_));
 sky130_fd_sc_hd__xnor2_1 _08446_ (.A(_01919_),
    .B(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__nand2_1 _08447_ (.A(_01801_),
    .B(_01804_),
    .Y(_01958_));
 sky130_fd_sc_hd__a21o_1 _08448_ (.A1(_01812_),
    .A2(_01820_),
    .B1(_01819_),
    .X(_01959_));
 sky130_fd_sc_hd__and4_1 _08449_ (.A(net36),
    .B(net37),
    .C(net11),
    .D(net13),
    .X(_01960_));
 sky130_fd_sc_hd__a22o_1 _08450_ (.A1(net37),
    .A2(net11),
    .B1(net13),
    .B2(net36),
    .X(_01961_));
 sky130_fd_sc_hd__and2b_1 _08451_ (.A_N(_01960_),
    .B(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__nand2_1 _08452_ (.A(net38),
    .B(net10),
    .Y(_01963_));
 sky130_fd_sc_hd__xnor2_1 _08453_ (.A(_01962_),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__nand4_1 _08454_ (.A(net64),
    .B(net34),
    .C(net15),
    .D(net16),
    .Y(_01965_));
 sky130_fd_sc_hd__a22o_1 _08455_ (.A1(net34),
    .A2(net15),
    .B1(net16),
    .B2(net64),
    .X(_01967_));
 sky130_fd_sc_hd__and2_1 _08456_ (.A(net35),
    .B(net14),
    .X(_01968_));
 sky130_fd_sc_hd__a21o_1 _08457_ (.A1(_01965_),
    .A2(_01967_),
    .B1(_01968_),
    .X(_01969_));
 sky130_fd_sc_hd__nand3_1 _08458_ (.A(_01965_),
    .B(_01967_),
    .C(_01968_),
    .Y(_01970_));
 sky130_fd_sc_hd__o21bai_1 _08459_ (.A1(_01622_),
    .A2(_01797_),
    .B1_N(_01796_),
    .Y(_01971_));
 sky130_fd_sc_hd__nand3_1 _08460_ (.A(_01969_),
    .B(_01970_),
    .C(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__a21o_1 _08461_ (.A1(_01969_),
    .A2(_01970_),
    .B1(_01971_),
    .X(_01973_));
 sky130_fd_sc_hd__nand3_1 _08462_ (.A(_01964_),
    .B(_01972_),
    .C(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__a21o_1 _08463_ (.A1(_01972_),
    .A2(_01973_),
    .B1(_01964_),
    .X(_01975_));
 sky130_fd_sc_hd__and3_1 _08464_ (.A(_01959_),
    .B(_01974_),
    .C(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__a21oi_1 _08465_ (.A1(_01974_),
    .A2(_01975_),
    .B1(_01959_),
    .Y(_01978_));
 sky130_fd_sc_hd__nor2_1 _08466_ (.A(_01976_),
    .B(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__xor2_1 _08467_ (.A(_01958_),
    .B(_01979_),
    .X(_01980_));
 sky130_fd_sc_hd__nand2_1 _08468_ (.A(_01816_),
    .B(_01818_),
    .Y(_01981_));
 sky130_fd_sc_hd__a22o_1 _08469_ (.A1(net21),
    .A2(_01823_),
    .B1(_01825_),
    .B2(_01652_),
    .X(_01982_));
 sky130_fd_sc_hd__nand4_1 _08470_ (.A(net61),
    .B(net62),
    .C(net18),
    .D(net19),
    .Y(_01983_));
 sky130_fd_sc_hd__a22o_1 _08471_ (.A1(net62),
    .A2(net18),
    .B1(net19),
    .B2(net61),
    .X(_01984_));
 sky130_fd_sc_hd__a22o_1 _08472_ (.A1(net63),
    .A2(net17),
    .B1(_01983_),
    .B2(_01984_),
    .X(_01985_));
 sky130_fd_sc_hd__nand4_1 _08473_ (.A(net63),
    .B(net17),
    .C(_01983_),
    .D(_01984_),
    .Y(_01986_));
 sky130_fd_sc_hd__and3_1 _08474_ (.A(_01982_),
    .B(_01985_),
    .C(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__a21o_1 _08475_ (.A1(_01985_),
    .A2(_01986_),
    .B1(_01982_),
    .X(_01989_));
 sky130_fd_sc_hd__and2b_1 _08476_ (.A_N(_01987_),
    .B(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__xor2_1 _08477_ (.A(_01981_),
    .B(_01990_),
    .X(_01991_));
 sky130_fd_sc_hd__nand2_1 _08478_ (.A(net60),
    .B(net20),
    .Y(_01992_));
 sky130_fd_sc_hd__and3_1 _08479_ (.A(net58),
    .B(net59),
    .C(net22),
    .X(_01993_));
 sky130_fd_sc_hd__and4_1 _08480_ (.A(net58),
    .B(net59),
    .C(net21),
    .D(net22),
    .X(_01994_));
 sky130_fd_sc_hd__a22o_1 _08481_ (.A1(net59),
    .A2(net21),
    .B1(net22),
    .B2(net58),
    .X(_01995_));
 sky130_fd_sc_hd__and2b_1 _08482_ (.A_N(_01994_),
    .B(_01995_),
    .X(_01996_));
 sky130_fd_sc_hd__xnor2_1 _08483_ (.A(_01992_),
    .B(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand3_2 _08484_ (.A(net33),
    .B(net44),
    .C(net25),
    .Y(_01998_));
 sky130_fd_sc_hd__o21a_1 _08485_ (.A1(net33),
    .A2(net44),
    .B1(net25),
    .X(_02000_));
 sky130_fd_sc_hd__o21ai_1 _08486_ (.A1(net33),
    .A2(net44),
    .B1(net25),
    .Y(_02001_));
 sky130_fd_sc_hd__a22o_1 _08487_ (.A1(net55),
    .A2(net24),
    .B1(_01998_),
    .B2(_02000_),
    .X(_02002_));
 sky130_fd_sc_hd__nand4_2 _08488_ (.A(net55),
    .B(net24),
    .C(_01998_),
    .D(_02000_),
    .Y(_02003_));
 sky130_fd_sc_hd__o21bai_1 _08489_ (.A1(_01658_),
    .A2(_01828_),
    .B1_N(_01829_),
    .Y(_02004_));
 sky130_fd_sc_hd__nand3_1 _08490_ (.A(_02002_),
    .B(_02003_),
    .C(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__a21o_1 _08491_ (.A1(_02002_),
    .A2(_02003_),
    .B1(_02004_),
    .X(_02006_));
 sky130_fd_sc_hd__nand3_1 _08492_ (.A(_01997_),
    .B(_02005_),
    .C(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__a21o_1 _08493_ (.A1(_02005_),
    .A2(_02006_),
    .B1(_01997_),
    .X(_02008_));
 sky130_fd_sc_hd__a21bo_1 _08494_ (.A1(_01827_),
    .A2(_01833_),
    .B1_N(_01832_),
    .X(_02009_));
 sky130_fd_sc_hd__nand3_1 _08495_ (.A(_02007_),
    .B(_02008_),
    .C(_02009_),
    .Y(_02011_));
 sky130_fd_sc_hd__a21o_1 _08496_ (.A1(_02007_),
    .A2(_02008_),
    .B1(_02009_),
    .X(_02012_));
 sky130_fd_sc_hd__and3_1 _08497_ (.A(_01991_),
    .B(_02011_),
    .C(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__a21oi_1 _08498_ (.A1(_02011_),
    .A2(_02012_),
    .B1(_01991_),
    .Y(_02014_));
 sky130_fd_sc_hd__a211o_1 _08499_ (.A1(_01838_),
    .A2(_01841_),
    .B1(_02013_),
    .C1(_02014_),
    .X(_02015_));
 sky130_fd_sc_hd__o211ai_2 _08500_ (.A1(_02013_),
    .A2(_02014_),
    .B1(_01838_),
    .C1(_01841_),
    .Y(_02016_));
 sky130_fd_sc_hd__nand3_1 _08501_ (.A(_01980_),
    .B(_02015_),
    .C(_02016_),
    .Y(_02017_));
 sky130_fd_sc_hd__a21o_1 _08502_ (.A1(_02015_),
    .A2(_02016_),
    .B1(_01980_),
    .X(_02018_));
 sky130_fd_sc_hd__o211a_1 _08503_ (.A1(_01843_),
    .A2(_01845_),
    .B1(_02017_),
    .C1(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__o211ai_1 _08504_ (.A1(_01843_),
    .A2(_01845_),
    .B1(_02017_),
    .C1(_02018_),
    .Y(_02020_));
 sky130_fd_sc_hd__a211o_1 _08505_ (.A1(_02017_),
    .A2(_02018_),
    .B1(_01843_),
    .C1(_01845_),
    .X(_02022_));
 sky130_fd_sc_hd__and3_1 _08506_ (.A(_01957_),
    .B(_02020_),
    .C(_02022_),
    .X(_02023_));
 sky130_fd_sc_hd__a21oi_1 _08507_ (.A1(_02020_),
    .A2(_02022_),
    .B1(_01957_),
    .Y(_02024_));
 sky130_fd_sc_hd__a211oi_1 _08508_ (.A1(_01848_),
    .A2(_01850_),
    .B1(_02023_),
    .C1(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__a211o_1 _08509_ (.A1(_01848_),
    .A2(_01850_),
    .B1(_02023_),
    .C1(_02024_),
    .X(_02026_));
 sky130_fd_sc_hd__o211ai_1 _08510_ (.A1(_02023_),
    .A2(_02024_),
    .B1(_01848_),
    .C1(_01850_),
    .Y(_02027_));
 sky130_fd_sc_hd__and3_1 _08511_ (.A(_01918_),
    .B(_02026_),
    .C(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__a21oi_1 _08512_ (.A1(_02026_),
    .A2(_02027_),
    .B1(_01918_),
    .Y(_02029_));
 sky130_fd_sc_hd__a211o_1 _08513_ (.A1(_01852_),
    .A2(_01854_),
    .B1(_02028_),
    .C1(_02029_),
    .X(_02030_));
 sky130_fd_sc_hd__o211ai_2 _08514_ (.A1(_02028_),
    .A2(_02029_),
    .B1(_01852_),
    .C1(_01854_),
    .Y(_02031_));
 sky130_fd_sc_hd__nand3_1 _08515_ (.A(_01871_),
    .B(_02030_),
    .C(_02031_),
    .Y(_02033_));
 sky130_fd_sc_hd__a21o_1 _08516_ (.A1(_02030_),
    .A2(_02031_),
    .B1(_01871_),
    .X(_02034_));
 sky130_fd_sc_hd__o211a_1 _08517_ (.A1(_01856_),
    .A2(_01859_),
    .B1(_02033_),
    .C1(_02034_),
    .X(_02035_));
 sky130_fd_sc_hd__o211ai_2 _08518_ (.A1(_01856_),
    .A2(_01859_),
    .B1(_02033_),
    .C1(_02034_),
    .Y(_02036_));
 sky130_fd_sc_hd__a211oi_1 _08519_ (.A1(_02033_),
    .A2(_02034_),
    .B1(_01856_),
    .C1(_01859_),
    .Y(_02037_));
 sky130_fd_sc_hd__or3_1 _08520_ (.A(_01724_),
    .B(_02035_),
    .C(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__o21ai_1 _08521_ (.A1(_02035_),
    .A2(_02037_),
    .B1(_01724_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand2_1 _08522_ (.A(_02038_),
    .B(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__and2b_1 _08523_ (.A_N(_01861_),
    .B(_01863_),
    .X(_02041_));
 sky130_fd_sc_hd__xnor2_1 _08524_ (.A(_02040_),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__or4bb_2 _08525_ (.A(_01867_),
    .B(_01702_),
    .C_N(_01699_),
    .D_N(_01866_),
    .X(_02044_));
 sky130_fd_sc_hd__and2_1 _08526_ (.A(_01065_),
    .B(_01218_),
    .X(_02045_));
 sky130_fd_sc_hd__a21o_1 _08527_ (.A1(_01698_),
    .A2(_01866_),
    .B1(_01867_),
    .X(_02046_));
 sky130_fd_sc_hd__a31o_1 _08528_ (.A1(_01699_),
    .A2(_01701_),
    .A3(_01869_),
    .B1(_02046_),
    .X(_02047_));
 sky130_fd_sc_hd__a21oi_2 _08529_ (.A1(_01067_),
    .A2(_02045_),
    .B1(_01220_),
    .Y(_02048_));
 sky130_fd_sc_hd__o21bai_4 _08530_ (.A1(_02044_),
    .A2(_02048_),
    .B1_N(_02047_),
    .Y(_02049_));
 sky130_fd_sc_hd__or3b_1 _08531_ (.A(_01068_),
    .B(_02044_),
    .C_N(_02045_),
    .X(_02050_));
 sky130_fd_sc_hd__and2b_2 _08532_ (.A_N(_02050_),
    .B(_00775_),
    .X(_02051_));
 sky130_fd_sc_hd__and3b_2 _08533_ (.A_N(_02050_),
    .B(_05524_),
    .C(_00776_),
    .X(_02052_));
 sky130_fd_sc_hd__or3_2 _08534_ (.A(_02049_),
    .B(_02051_),
    .C(_02052_),
    .X(_02053_));
 sky130_fd_sc_hd__nand2b_1 _08535_ (.A_N(_02042_),
    .B(_02053_),
    .Y(_02055_));
 sky130_fd_sc_hd__xnor2_1 _08536_ (.A(_02042_),
    .B(_02053_),
    .Y(net90));
 sky130_fd_sc_hd__nand2_1 _08537_ (.A(_01890_),
    .B(_01892_),
    .Y(_02056_));
 sky130_fd_sc_hd__a21o_1 _08538_ (.A1(_01872_),
    .A2(_01917_),
    .B1(_01916_),
    .X(_02057_));
 sky130_fd_sc_hd__o21ba_1 _08539_ (.A1(_01894_),
    .A2(_01913_),
    .B1_N(_01912_),
    .X(_02058_));
 sky130_fd_sc_hd__o21ba_1 _08540_ (.A1(_01919_),
    .A2(_01954_),
    .B1_N(_01953_),
    .X(_02059_));
 sky130_fd_sc_hd__and4_1 _08541_ (.A(net28),
    .B(net29),
    .C(net52),
    .D(net53),
    .X(_02060_));
 sky130_fd_sc_hd__a22oi_1 _08542_ (.A1(net29),
    .A2(net52),
    .B1(net53),
    .B2(net28),
    .Y(_02061_));
 sky130_fd_sc_hd__nor2_1 _08543_ (.A(_02060_),
    .B(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__nand2_1 _08544_ (.A(net27),
    .B(net54),
    .Y(_02063_));
 sky130_fd_sc_hd__xnor2_1 _08545_ (.A(_02062_),
    .B(_02063_),
    .Y(_02065_));
 sky130_fd_sc_hd__a31o_1 _08546_ (.A1(net26),
    .A2(net54),
    .A3(_01880_),
    .B1(_01879_),
    .X(_02066_));
 sky130_fd_sc_hd__and2_1 _08547_ (.A(_02065_),
    .B(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__xor2_1 _08548_ (.A(_02065_),
    .B(_02066_),
    .X(_02068_));
 sky130_fd_sc_hd__and4b_1 _08549_ (.A_N(net23),
    .B(net56),
    .C(net57),
    .D(net26),
    .X(_02069_));
 sky130_fd_sc_hd__inv_2 _08550_ (.A(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__o2bb2a_1 _08551_ (.A1_N(net26),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net23),
    .X(_02071_));
 sky130_fd_sc_hd__nor2_1 _08552_ (.A(_02069_),
    .B(_02071_),
    .Y(_02072_));
 sky130_fd_sc_hd__xnor2_1 _08553_ (.A(_02068_),
    .B(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__and3_1 _08554_ (.A(_01885_),
    .B(_01887_),
    .C(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__a21o_1 _08555_ (.A1(_01885_),
    .A2(_01887_),
    .B1(_02073_),
    .X(_02076_));
 sky130_fd_sc_hd__nand2b_1 _08556_ (.A_N(_02074_),
    .B(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__xnor2_1 _08557_ (.A(_01875_),
    .B(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__a21o_1 _08558_ (.A1(_01925_),
    .A2(_01934_),
    .B1(_01932_),
    .X(_02079_));
 sky130_fd_sc_hd__nand2_1 _08559_ (.A(_01898_),
    .B(_01902_),
    .Y(_02080_));
 sky130_fd_sc_hd__a31o_1 _08560_ (.A1(net32),
    .A2(net48),
    .A3(_01921_),
    .B1(_01920_),
    .X(_02081_));
 sky130_fd_sc_hd__nand4_1 _08561_ (.A(net31),
    .B(net32),
    .C(net49),
    .D(net50),
    .Y(_02082_));
 sky130_fd_sc_hd__a22o_1 _08562_ (.A1(net32),
    .A2(net49),
    .B1(net50),
    .B2(net31),
    .X(_02083_));
 sky130_fd_sc_hd__a22o_1 _08563_ (.A1(net30),
    .A2(net51),
    .B1(_02082_),
    .B2(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__nand4_1 _08564_ (.A(net30),
    .B(net51),
    .C(_02082_),
    .D(_02083_),
    .Y(_02085_));
 sky130_fd_sc_hd__nand3_1 _08565_ (.A(_02081_),
    .B(_02084_),
    .C(_02085_),
    .Y(_02087_));
 sky130_fd_sc_hd__a21o_1 _08566_ (.A1(_02084_),
    .A2(_02085_),
    .B1(_02081_),
    .X(_02088_));
 sky130_fd_sc_hd__nand3_1 _08567_ (.A(_02080_),
    .B(_02087_),
    .C(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__a21o_1 _08568_ (.A1(_02087_),
    .A2(_02088_),
    .B1(_02080_),
    .X(_02090_));
 sky130_fd_sc_hd__and3_1 _08569_ (.A(_02079_),
    .B(_02089_),
    .C(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__a21oi_1 _08570_ (.A1(_02089_),
    .A2(_02090_),
    .B1(_02079_),
    .Y(_02092_));
 sky130_fd_sc_hd__a211oi_1 _08571_ (.A1(_01903_),
    .A2(_01905_),
    .B1(_02091_),
    .C1(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__o211a_1 _08572_ (.A1(_02091_),
    .A2(_02092_),
    .B1(_01903_),
    .C1(_01905_),
    .X(_02094_));
 sky130_fd_sc_hd__or2_1 _08573_ (.A(_02093_),
    .B(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__and2b_1 _08574_ (.A_N(_01907_),
    .B(_01909_),
    .X(_02096_));
 sky130_fd_sc_hd__nor2_1 _08575_ (.A(_02095_),
    .B(_02096_),
    .Y(_02098_));
 sky130_fd_sc_hd__xnor2_1 _08576_ (.A(_02095_),
    .B(_02096_),
    .Y(_02099_));
 sky130_fd_sc_hd__xnor2_1 _08577_ (.A(_02078_),
    .B(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__xor2_1 _08578_ (.A(_02059_),
    .B(_02100_),
    .X(_02101_));
 sky130_fd_sc_hd__nand2b_1 _08579_ (.A_N(_02058_),
    .B(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hd__xnor2_1 _08580_ (.A(_02058_),
    .B(_02101_),
    .Y(_02103_));
 sky130_fd_sc_hd__or2_1 _08581_ (.A(_01949_),
    .B(_01951_),
    .X(_02104_));
 sky130_fd_sc_hd__a21oi_1 _08582_ (.A1(_01958_),
    .A2(_01979_),
    .B1(_01976_),
    .Y(_02105_));
 sky130_fd_sc_hd__and4_1 _08583_ (.A(net3),
    .B(net4),
    .C(net46),
    .D(net47),
    .X(_02106_));
 sky130_fd_sc_hd__a22o_1 _08584_ (.A1(net4),
    .A2(net46),
    .B1(net47),
    .B2(net3),
    .X(_02107_));
 sky130_fd_sc_hd__and2b_1 _08585_ (.A_N(_02106_),
    .B(_02107_),
    .X(_02109_));
 sky130_fd_sc_hd__nand2_1 _08586_ (.A(net2),
    .B(net48),
    .Y(_02110_));
 sky130_fd_sc_hd__xnor2_1 _08587_ (.A(_02109_),
    .B(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__nand2_1 _08588_ (.A(net5),
    .B(net45),
    .Y(_02112_));
 sky130_fd_sc_hd__and4_1 _08589_ (.A(net6),
    .B(net7),
    .C(net42),
    .D(net43),
    .X(_02113_));
 sky130_fd_sc_hd__a22oi_2 _08590_ (.A1(net7),
    .A2(net42),
    .B1(net43),
    .B2(net6),
    .Y(_02114_));
 sky130_fd_sc_hd__or3_1 _08591_ (.A(_02112_),
    .B(_02113_),
    .C(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__o21ai_1 _08592_ (.A1(_02113_),
    .A2(_02114_),
    .B1(_02112_),
    .Y(_02116_));
 sky130_fd_sc_hd__a21bo_1 _08593_ (.A1(_01927_),
    .A2(_01928_),
    .B1_N(_01926_),
    .X(_02117_));
 sky130_fd_sc_hd__and3_1 _08594_ (.A(_02115_),
    .B(_02116_),
    .C(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__a21o_1 _08595_ (.A1(_02115_),
    .A2(_02116_),
    .B1(_02117_),
    .X(_02120_));
 sky130_fd_sc_hd__and2b_1 _08596_ (.A_N(_02118_),
    .B(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__xnor2_1 _08597_ (.A(_02111_),
    .B(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_1 _08598_ (.A(_01939_),
    .B(_01942_),
    .Y(_02123_));
 sky130_fd_sc_hd__a31o_1 _08599_ (.A1(net38),
    .A2(net10),
    .A3(_01961_),
    .B1(_01960_),
    .X(_02124_));
 sky130_fd_sc_hd__nand4_1 _08600_ (.A(net39),
    .B(net40),
    .C(net9),
    .D(net10),
    .Y(_02125_));
 sky130_fd_sc_hd__a22o_1 _08601_ (.A1(net40),
    .A2(net9),
    .B1(net10),
    .B2(net39),
    .X(_02126_));
 sky130_fd_sc_hd__a22o_1 _08602_ (.A1(net8),
    .A2(net41),
    .B1(_02125_),
    .B2(_02126_),
    .X(_02127_));
 sky130_fd_sc_hd__nand4_1 _08603_ (.A(net8),
    .B(net41),
    .C(_02125_),
    .D(_02126_),
    .Y(_02128_));
 sky130_fd_sc_hd__nand3_1 _08604_ (.A(_02124_),
    .B(_02127_),
    .C(_02128_),
    .Y(_02129_));
 sky130_fd_sc_hd__a21o_1 _08605_ (.A1(_02127_),
    .A2(_02128_),
    .B1(_02124_),
    .X(_02131_));
 sky130_fd_sc_hd__nand3_1 _08606_ (.A(_02123_),
    .B(_02129_),
    .C(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__a21o_1 _08607_ (.A1(_02129_),
    .A2(_02131_),
    .B1(_02123_),
    .X(_02133_));
 sky130_fd_sc_hd__a21bo_1 _08608_ (.A1(_01937_),
    .A2(_01945_),
    .B1_N(_01943_),
    .X(_02134_));
 sky130_fd_sc_hd__and3_1 _08609_ (.A(_02132_),
    .B(_02133_),
    .C(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__a21oi_1 _08610_ (.A1(_02132_),
    .A2(_02133_),
    .B1(_02134_),
    .Y(_02136_));
 sky130_fd_sc_hd__nor3_1 _08611_ (.A(_02122_),
    .B(_02135_),
    .C(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__o21a_1 _08612_ (.A1(_02135_),
    .A2(_02136_),
    .B1(_02122_),
    .X(_02138_));
 sky130_fd_sc_hd__or2_1 _08613_ (.A(_02137_),
    .B(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__or2_1 _08614_ (.A(_02105_),
    .B(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__xor2_1 _08615_ (.A(_02105_),
    .B(_02139_),
    .X(_02142_));
 sky130_fd_sc_hd__xor2_1 _08616_ (.A(_02104_),
    .B(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__nand2_1 _08617_ (.A(_01972_),
    .B(_01974_),
    .Y(_02144_));
 sky130_fd_sc_hd__a21o_1 _08618_ (.A1(_01981_),
    .A2(_01989_),
    .B1(_01987_),
    .X(_02145_));
 sky130_fd_sc_hd__nand2_1 _08619_ (.A(net38),
    .B(net11),
    .Y(_02146_));
 sky130_fd_sc_hd__and4_1 _08620_ (.A(net36),
    .B(net37),
    .C(net13),
    .D(net14),
    .X(_02147_));
 sky130_fd_sc_hd__a22o_1 _08621_ (.A1(net37),
    .A2(net13),
    .B1(net14),
    .B2(net36),
    .X(_02148_));
 sky130_fd_sc_hd__and2b_1 _08622_ (.A_N(_02147_),
    .B(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__xnor2_1 _08623_ (.A(_02146_),
    .B(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__nand2_1 _08624_ (.A(net35),
    .B(net15),
    .Y(_02151_));
 sky130_fd_sc_hd__and4_1 _08625_ (.A(net64),
    .B(net34),
    .C(net16),
    .D(net17),
    .X(_02153_));
 sky130_fd_sc_hd__a22oi_2 _08626_ (.A1(net34),
    .A2(net16),
    .B1(net17),
    .B2(net64),
    .Y(_02154_));
 sky130_fd_sc_hd__or3_1 _08627_ (.A(_02151_),
    .B(_02153_),
    .C(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__o21ai_1 _08628_ (.A1(_02153_),
    .A2(_02154_),
    .B1(_02151_),
    .Y(_02156_));
 sky130_fd_sc_hd__a21bo_1 _08629_ (.A1(_01967_),
    .A2(_01968_),
    .B1_N(_01965_),
    .X(_02157_));
 sky130_fd_sc_hd__nand3_2 _08630_ (.A(_02155_),
    .B(_02156_),
    .C(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__a21o_1 _08631_ (.A1(_02155_),
    .A2(_02156_),
    .B1(_02157_),
    .X(_02159_));
 sky130_fd_sc_hd__nand3_1 _08632_ (.A(_02150_),
    .B(_02158_),
    .C(_02159_),
    .Y(_02160_));
 sky130_fd_sc_hd__a21o_1 _08633_ (.A1(_02158_),
    .A2(_02159_),
    .B1(_02150_),
    .X(_02161_));
 sky130_fd_sc_hd__and3_1 _08634_ (.A(_02145_),
    .B(_02160_),
    .C(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__a21oi_1 _08635_ (.A1(_02160_),
    .A2(_02161_),
    .B1(_02145_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_1 _08636_ (.A(_02162_),
    .B(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__xor2_1 _08637_ (.A(_02144_),
    .B(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__nand2_1 _08638_ (.A(_01983_),
    .B(_01986_),
    .Y(_02167_));
 sky130_fd_sc_hd__a31o_1 _08639_ (.A1(net60),
    .A2(net20),
    .A3(_01995_),
    .B1(_01994_),
    .X(_02168_));
 sky130_fd_sc_hd__nand2_1 _08640_ (.A(net63),
    .B(net18),
    .Y(_02169_));
 sky130_fd_sc_hd__nand4_1 _08641_ (.A(net61),
    .B(net62),
    .C(net19),
    .D(net20),
    .Y(_02170_));
 sky130_fd_sc_hd__a22o_1 _08642_ (.A1(net62),
    .A2(net19),
    .B1(net20),
    .B2(net61),
    .X(_02171_));
 sky130_fd_sc_hd__nand3b_1 _08643_ (.A_N(_02169_),
    .B(_02170_),
    .C(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__a21bo_1 _08644_ (.A1(_02170_),
    .A2(_02171_),
    .B1_N(_02169_),
    .X(_02173_));
 sky130_fd_sc_hd__and3_1 _08645_ (.A(_02168_),
    .B(_02172_),
    .C(_02173_),
    .X(_02175_));
 sky130_fd_sc_hd__a21o_1 _08646_ (.A1(_02172_),
    .A2(_02173_),
    .B1(_02168_),
    .X(_02176_));
 sky130_fd_sc_hd__and2b_1 _08647_ (.A_N(_02175_),
    .B(_02176_),
    .X(_02177_));
 sky130_fd_sc_hd__xnor2_1 _08648_ (.A(_02167_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__nand2_1 _08649_ (.A(net60),
    .B(net21),
    .Y(_02179_));
 sky130_fd_sc_hd__a22o_1 _08650_ (.A1(net59),
    .A2(net22),
    .B1(net24),
    .B2(net58),
    .X(_02180_));
 sky130_fd_sc_hd__a21bo_1 _08651_ (.A1(net24),
    .A2(_01993_),
    .B1_N(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__xor2_1 _08652_ (.A(_02179_),
    .B(_02181_),
    .X(_02182_));
 sky130_fd_sc_hd__nand2_1 _08653_ (.A(net55),
    .B(net25),
    .Y(_02183_));
 sky130_fd_sc_hd__nand3_1 _08654_ (.A(_01998_),
    .B(_02000_),
    .C(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__a21o_1 _08655_ (.A1(_01998_),
    .A2(_02000_),
    .B1(_02183_),
    .X(_02186_));
 sky130_fd_sc_hd__nand4_1 _08656_ (.A(_01998_),
    .B(_02003_),
    .C(_02184_),
    .D(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__and4_2 _08657_ (.A(net33),
    .B(net44),
    .C(net55),
    .D(net25),
    .X(_02188_));
 sky130_fd_sc_hd__a41o_1 _08658_ (.A1(_01998_),
    .A2(_02003_),
    .A3(_02184_),
    .A4(_02186_),
    .B1(_02188_),
    .X(_02189_));
 sky130_fd_sc_hd__xor2_1 _08659_ (.A(_02182_),
    .B(_02189_),
    .X(_02190_));
 sky130_fd_sc_hd__a21bo_1 _08660_ (.A1(_01997_),
    .A2(_02006_),
    .B1_N(_02005_),
    .X(_02191_));
 sky130_fd_sc_hd__nand2b_1 _08661_ (.A_N(_02190_),
    .B(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__xor2_1 _08662_ (.A(_02190_),
    .B(_02191_),
    .X(_02193_));
 sky130_fd_sc_hd__xnor2_1 _08663_ (.A(_02178_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__a21boi_1 _08664_ (.A1(_01991_),
    .A2(_02012_),
    .B1_N(_02011_),
    .Y(_02195_));
 sky130_fd_sc_hd__nor2_1 _08665_ (.A(_02194_),
    .B(_02195_),
    .Y(_02197_));
 sky130_fd_sc_hd__xor2_1 _08666_ (.A(_02194_),
    .B(_02195_),
    .X(_02198_));
 sky130_fd_sc_hd__xnor2_1 _08667_ (.A(_02166_),
    .B(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__a21bo_1 _08668_ (.A1(_01980_),
    .A2(_02016_),
    .B1_N(_02015_),
    .X(_02200_));
 sky130_fd_sc_hd__and2b_1 _08669_ (.A_N(_02199_),
    .B(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__xnor2_1 _08670_ (.A(_02199_),
    .B(_02200_),
    .Y(_02202_));
 sky130_fd_sc_hd__xor2_1 _08671_ (.A(_02143_),
    .B(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__a21oi_1 _08672_ (.A1(_01957_),
    .A2(_02022_),
    .B1(_02019_),
    .Y(_02204_));
 sky130_fd_sc_hd__and2b_1 _08673_ (.A_N(_02204_),
    .B(_02203_),
    .X(_02205_));
 sky130_fd_sc_hd__xnor2_1 _08674_ (.A(_02203_),
    .B(_02204_),
    .Y(_02206_));
 sky130_fd_sc_hd__xor2_1 _08675_ (.A(_02103_),
    .B(_02206_),
    .X(_02207_));
 sky130_fd_sc_hd__a21oi_1 _08676_ (.A1(_01918_),
    .A2(_02027_),
    .B1(_02025_),
    .Y(_02208_));
 sky130_fd_sc_hd__and2b_1 _08677_ (.A_N(_02208_),
    .B(_02207_),
    .X(_02209_));
 sky130_fd_sc_hd__xnor2_1 _08678_ (.A(_02207_),
    .B(_02208_),
    .Y(_02210_));
 sky130_fd_sc_hd__xnor2_2 _08679_ (.A(_02057_),
    .B(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__a21boi_2 _08680_ (.A1(_01871_),
    .A2(_02031_),
    .B1_N(_02030_),
    .Y(_02212_));
 sky130_fd_sc_hd__nor2_1 _08681_ (.A(_02211_),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__xor2_2 _08682_ (.A(_02211_),
    .B(_02212_),
    .X(_02214_));
 sky130_fd_sc_hd__xnor2_1 _08683_ (.A(_02056_),
    .B(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__a21oi_1 _08684_ (.A1(_02036_),
    .A2(_02038_),
    .B1(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__a21o_1 _08685_ (.A1(_02036_),
    .A2(_02038_),
    .B1(_02215_),
    .X(_02218_));
 sky130_fd_sc_hd__and3_1 _08686_ (.A(_02036_),
    .B(_02038_),
    .C(_02215_),
    .X(_02219_));
 sky130_fd_sc_hd__or2_1 _08687_ (.A(_02216_),
    .B(_02219_),
    .X(_02220_));
 sky130_fd_sc_hd__o21ai_1 _08688_ (.A1(_02040_),
    .A2(_02041_),
    .B1(_02055_),
    .Y(_02221_));
 sky130_fd_sc_hd__xnor2_1 _08689_ (.A(_02220_),
    .B(_02221_),
    .Y(net91));
 sky130_fd_sc_hd__o21ai_1 _08690_ (.A1(_01875_),
    .A2(_02074_),
    .B1(_02076_),
    .Y(_02222_));
 sky130_fd_sc_hd__o21ai_1 _08691_ (.A1(_02059_),
    .A2(_02100_),
    .B1(_02102_),
    .Y(_02223_));
 sky130_fd_sc_hd__o21ba_1 _08692_ (.A1(_02078_),
    .A2(_02099_),
    .B1_N(_02098_),
    .X(_02224_));
 sky130_fd_sc_hd__a21boi_1 _08693_ (.A1(_02104_),
    .A2(_02142_),
    .B1_N(_02140_),
    .Y(_02225_));
 sky130_fd_sc_hd__and4_1 _08694_ (.A(net29),
    .B(net30),
    .C(net52),
    .D(net53),
    .X(_02226_));
 sky130_fd_sc_hd__a22oi_1 _08695_ (.A1(net30),
    .A2(net52),
    .B1(net53),
    .B2(net29),
    .Y(_02228_));
 sky130_fd_sc_hd__nor2_1 _08696_ (.A(_02226_),
    .B(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__nand2_1 _08697_ (.A(net28),
    .B(net54),
    .Y(_02230_));
 sky130_fd_sc_hd__xnor2_1 _08698_ (.A(_02229_),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__o21ba_1 _08699_ (.A1(_02061_),
    .A2(_02063_),
    .B1_N(_02060_),
    .X(_02232_));
 sky130_fd_sc_hd__nand2b_1 _08700_ (.A_N(_02232_),
    .B(_02231_),
    .Y(_02233_));
 sky130_fd_sc_hd__xnor2_1 _08701_ (.A(_02231_),
    .B(_02232_),
    .Y(_02234_));
 sky130_fd_sc_hd__and4b_1 _08702_ (.A_N(net26),
    .B(net56),
    .C(net57),
    .D(net27),
    .X(_02235_));
 sky130_fd_sc_hd__inv_2 _08703_ (.A(_02235_),
    .Y(_02236_));
 sky130_fd_sc_hd__o2bb2a_1 _08704_ (.A1_N(net27),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net26),
    .X(_02237_));
 sky130_fd_sc_hd__nor2_1 _08705_ (.A(_02235_),
    .B(_02237_),
    .Y(_02239_));
 sky130_fd_sc_hd__or2_1 _08706_ (.A(_02234_),
    .B(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__nand2_1 _08707_ (.A(_02234_),
    .B(_02239_),
    .Y(_02241_));
 sky130_fd_sc_hd__nand2_1 _08708_ (.A(_02240_),
    .B(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__a21o_1 _08709_ (.A1(_02068_),
    .A2(_02072_),
    .B1(_02067_),
    .X(_02243_));
 sky130_fd_sc_hd__nand2b_1 _08710_ (.A_N(_02242_),
    .B(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__xor2_1 _08711_ (.A(_02242_),
    .B(_02243_),
    .X(_02245_));
 sky130_fd_sc_hd__xnor2_1 _08712_ (.A(_02070_),
    .B(_02245_),
    .Y(_02246_));
 sky130_fd_sc_hd__a21o_1 _08713_ (.A1(_02111_),
    .A2(_02120_),
    .B1(_02118_),
    .X(_02247_));
 sky130_fd_sc_hd__nand2_1 _08714_ (.A(_02082_),
    .B(_02085_),
    .Y(_02248_));
 sky130_fd_sc_hd__a31o_1 _08715_ (.A1(net2),
    .A2(net48),
    .A3(_02107_),
    .B1(_02106_),
    .X(_02250_));
 sky130_fd_sc_hd__nand4_1 _08716_ (.A(net2),
    .B(net32),
    .C(net49),
    .D(net50),
    .Y(_02251_));
 sky130_fd_sc_hd__a22o_1 _08717_ (.A1(net2),
    .A2(net49),
    .B1(net50),
    .B2(net32),
    .X(_02252_));
 sky130_fd_sc_hd__a22o_1 _08718_ (.A1(net31),
    .A2(net51),
    .B1(_02251_),
    .B2(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__nand4_1 _08719_ (.A(net31),
    .B(net51),
    .C(_02251_),
    .D(_02252_),
    .Y(_02254_));
 sky130_fd_sc_hd__nand3_1 _08720_ (.A(_02250_),
    .B(_02253_),
    .C(_02254_),
    .Y(_02255_));
 sky130_fd_sc_hd__a21o_1 _08721_ (.A1(_02253_),
    .A2(_02254_),
    .B1(_02250_),
    .X(_02256_));
 sky130_fd_sc_hd__nand3_1 _08722_ (.A(_02248_),
    .B(_02255_),
    .C(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__a21o_1 _08723_ (.A1(_02255_),
    .A2(_02256_),
    .B1(_02248_),
    .X(_02258_));
 sky130_fd_sc_hd__and3_1 _08724_ (.A(_02247_),
    .B(_02257_),
    .C(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__a21oi_1 _08725_ (.A1(_02257_),
    .A2(_02258_),
    .B1(_02247_),
    .Y(_02261_));
 sky130_fd_sc_hd__a211oi_1 _08726_ (.A1(_02087_),
    .A2(_02089_),
    .B1(_02259_),
    .C1(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__o211a_1 _08727_ (.A1(_02259_),
    .A2(_02261_),
    .B1(_02087_),
    .C1(_02089_),
    .X(_02263_));
 sky130_fd_sc_hd__or2_1 _08728_ (.A(_02262_),
    .B(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__nor2_1 _08729_ (.A(_02091_),
    .B(_02093_),
    .Y(_02265_));
 sky130_fd_sc_hd__nor2_1 _08730_ (.A(_02264_),
    .B(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__xnor2_1 _08731_ (.A(_02264_),
    .B(_02265_),
    .Y(_02267_));
 sky130_fd_sc_hd__xnor2_1 _08732_ (.A(_02246_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__xor2_1 _08733_ (.A(_02225_),
    .B(_02268_),
    .X(_02269_));
 sky130_fd_sc_hd__and2b_1 _08734_ (.A_N(_02224_),
    .B(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__xnor2_1 _08735_ (.A(_02224_),
    .B(_02269_),
    .Y(_02272_));
 sky130_fd_sc_hd__or2_1 _08736_ (.A(_02135_),
    .B(_02137_),
    .X(_02273_));
 sky130_fd_sc_hd__a21o_1 _08737_ (.A1(_02144_),
    .A2(_02165_),
    .B1(_02162_),
    .X(_02274_));
 sky130_fd_sc_hd__and4_1 _08738_ (.A(net4),
    .B(net5),
    .C(net46),
    .D(net47),
    .X(_02275_));
 sky130_fd_sc_hd__a22o_1 _08739_ (.A1(net5),
    .A2(net46),
    .B1(net47),
    .B2(net4),
    .X(_02276_));
 sky130_fd_sc_hd__and2b_1 _08740_ (.A_N(_02275_),
    .B(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__nand2_1 _08741_ (.A(net3),
    .B(net48),
    .Y(_02278_));
 sky130_fd_sc_hd__xnor2_1 _08742_ (.A(_02277_),
    .B(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__nand2_1 _08743_ (.A(net6),
    .B(net45),
    .Y(_02280_));
 sky130_fd_sc_hd__and4_1 _08744_ (.A(net7),
    .B(net8),
    .C(net42),
    .D(net43),
    .X(_02281_));
 sky130_fd_sc_hd__a22oi_2 _08745_ (.A1(net8),
    .A2(net42),
    .B1(net43),
    .B2(net7),
    .Y(_02283_));
 sky130_fd_sc_hd__or3_1 _08746_ (.A(_02280_),
    .B(_02281_),
    .C(_02283_),
    .X(_02284_));
 sky130_fd_sc_hd__o21ai_1 _08747_ (.A1(_02281_),
    .A2(_02283_),
    .B1(_02280_),
    .Y(_02285_));
 sky130_fd_sc_hd__o21bai_1 _08748_ (.A1(_02112_),
    .A2(_02114_),
    .B1_N(_02113_),
    .Y(_02286_));
 sky130_fd_sc_hd__and3_1 _08749_ (.A(_02284_),
    .B(_02285_),
    .C(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__a21o_1 _08750_ (.A1(_02284_),
    .A2(_02285_),
    .B1(_02286_),
    .X(_02288_));
 sky130_fd_sc_hd__and2b_1 _08751_ (.A_N(_02287_),
    .B(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__xnor2_1 _08752_ (.A(_02279_),
    .B(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__nand2_1 _08753_ (.A(_02125_),
    .B(_02128_),
    .Y(_02291_));
 sky130_fd_sc_hd__a31o_1 _08754_ (.A1(net38),
    .A2(net11),
    .A3(_02148_),
    .B1(_02147_),
    .X(_02292_));
 sky130_fd_sc_hd__nand4_1 _08755_ (.A(net39),
    .B(net40),
    .C(net10),
    .D(net11),
    .Y(_02294_));
 sky130_fd_sc_hd__a22o_1 _08756_ (.A1(net40),
    .A2(net10),
    .B1(net11),
    .B2(net39),
    .X(_02295_));
 sky130_fd_sc_hd__a22o_1 _08757_ (.A1(net9),
    .A2(net41),
    .B1(_02294_),
    .B2(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__nand4_1 _08758_ (.A(net9),
    .B(net41),
    .C(_02294_),
    .D(_02295_),
    .Y(_02297_));
 sky130_fd_sc_hd__nand3_1 _08759_ (.A(_02292_),
    .B(_02296_),
    .C(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__a21o_1 _08760_ (.A1(_02296_),
    .A2(_02297_),
    .B1(_02292_),
    .X(_02299_));
 sky130_fd_sc_hd__nand3_1 _08761_ (.A(_02291_),
    .B(_02298_),
    .C(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__a21o_1 _08762_ (.A1(_02298_),
    .A2(_02299_),
    .B1(_02291_),
    .X(_02301_));
 sky130_fd_sc_hd__a21bo_1 _08763_ (.A1(_02123_),
    .A2(_02131_),
    .B1_N(_02129_),
    .X(_02302_));
 sky130_fd_sc_hd__and3_1 _08764_ (.A(_02300_),
    .B(_02301_),
    .C(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__a21oi_1 _08765_ (.A1(_02300_),
    .A2(_02301_),
    .B1(_02302_),
    .Y(_02305_));
 sky130_fd_sc_hd__nor3_1 _08766_ (.A(_02290_),
    .B(_02303_),
    .C(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__o21a_1 _08767_ (.A1(_02303_),
    .A2(_02305_),
    .B1(_02290_),
    .X(_02307_));
 sky130_fd_sc_hd__or2_1 _08768_ (.A(_02306_),
    .B(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__nand2b_1 _08769_ (.A_N(_02308_),
    .B(_02274_),
    .Y(_02309_));
 sky130_fd_sc_hd__xnor2_1 _08770_ (.A(_02274_),
    .B(_02308_),
    .Y(_02310_));
 sky130_fd_sc_hd__xor2_1 _08771_ (.A(_02273_),
    .B(_02310_),
    .X(_02311_));
 sky130_fd_sc_hd__a21o_1 _08772_ (.A1(_02167_),
    .A2(_02176_),
    .B1(_02175_),
    .X(_02312_));
 sky130_fd_sc_hd__nand2_1 _08773_ (.A(net38),
    .B(net13),
    .Y(_02313_));
 sky130_fd_sc_hd__and4_1 _08774_ (.A(net36),
    .B(net37),
    .C(net14),
    .D(net15),
    .X(_02314_));
 sky130_fd_sc_hd__a22o_1 _08775_ (.A1(net37),
    .A2(net14),
    .B1(net15),
    .B2(net36),
    .X(_02316_));
 sky130_fd_sc_hd__and2b_1 _08776_ (.A_N(_02314_),
    .B(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__xnor2_1 _08777_ (.A(_02313_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__nand2_1 _08778_ (.A(net35),
    .B(net16),
    .Y(_02319_));
 sky130_fd_sc_hd__and4_1 _08779_ (.A(net64),
    .B(net34),
    .C(net17),
    .D(net18),
    .X(_02320_));
 sky130_fd_sc_hd__a22oi_2 _08780_ (.A1(net34),
    .A2(net17),
    .B1(net18),
    .B2(net64),
    .Y(_02321_));
 sky130_fd_sc_hd__or3_1 _08781_ (.A(_02319_),
    .B(_02320_),
    .C(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__o21ai_1 _08782_ (.A1(_02320_),
    .A2(_02321_),
    .B1(_02319_),
    .Y(_02323_));
 sky130_fd_sc_hd__o21bai_1 _08783_ (.A1(_02151_),
    .A2(_02154_),
    .B1_N(_02153_),
    .Y(_02324_));
 sky130_fd_sc_hd__nand3_1 _08784_ (.A(_02322_),
    .B(_02323_),
    .C(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__a21o_1 _08785_ (.A1(_02322_),
    .A2(_02323_),
    .B1(_02324_),
    .X(_02327_));
 sky130_fd_sc_hd__nand3_1 _08786_ (.A(_02318_),
    .B(_02325_),
    .C(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__a21o_1 _08787_ (.A1(_02325_),
    .A2(_02327_),
    .B1(_02318_),
    .X(_02329_));
 sky130_fd_sc_hd__and3_1 _08788_ (.A(_02312_),
    .B(_02328_),
    .C(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__a21oi_1 _08789_ (.A1(_02328_),
    .A2(_02329_),
    .B1(_02312_),
    .Y(_02331_));
 sky130_fd_sc_hd__a211oi_2 _08790_ (.A1(_02158_),
    .A2(_02160_),
    .B1(_02330_),
    .C1(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__o211a_1 _08791_ (.A1(_02330_),
    .A2(_02331_),
    .B1(_02158_),
    .C1(_02160_),
    .X(_02333_));
 sky130_fd_sc_hd__nor2_1 _08792_ (.A(_02332_),
    .B(_02333_),
    .Y(_02334_));
 sky130_fd_sc_hd__nand2_1 _08793_ (.A(_02170_),
    .B(_02172_),
    .Y(_02335_));
 sky130_fd_sc_hd__a32o_1 _08794_ (.A1(net60),
    .A2(net21),
    .A3(_02180_),
    .B1(_01993_),
    .B2(net24),
    .X(_02336_));
 sky130_fd_sc_hd__nand2_1 _08795_ (.A(net63),
    .B(net19),
    .Y(_02338_));
 sky130_fd_sc_hd__nand4_1 _08796_ (.A(net61),
    .B(net62),
    .C(net20),
    .D(net21),
    .Y(_02339_));
 sky130_fd_sc_hd__a22o_1 _08797_ (.A1(net62),
    .A2(net20),
    .B1(net21),
    .B2(net61),
    .X(_02340_));
 sky130_fd_sc_hd__nand3b_1 _08798_ (.A_N(_02338_),
    .B(_02339_),
    .C(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__a21bo_1 _08799_ (.A1(_02339_),
    .A2(_02340_),
    .B1_N(_02338_),
    .X(_02342_));
 sky130_fd_sc_hd__and3_1 _08800_ (.A(_02336_),
    .B(_02341_),
    .C(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__a21o_1 _08801_ (.A1(_02341_),
    .A2(_02342_),
    .B1(_02336_),
    .X(_02344_));
 sky130_fd_sc_hd__and2b_1 _08802_ (.A_N(_02343_),
    .B(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__xnor2_1 _08803_ (.A(_02335_),
    .B(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__nand2_1 _08804_ (.A(net60),
    .B(net22),
    .Y(_02347_));
 sky130_fd_sc_hd__and4_1 _08805_ (.A(net58),
    .B(net59),
    .C(net24),
    .D(net25),
    .X(_02349_));
 sky130_fd_sc_hd__a22oi_2 _08806_ (.A1(net59),
    .A2(net24),
    .B1(net25),
    .B2(net58),
    .Y(_02350_));
 sky130_fd_sc_hd__or3_1 _08807_ (.A(_02347_),
    .B(_02349_),
    .C(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__o21ai_1 _08808_ (.A1(_02349_),
    .A2(_02350_),
    .B1(_02347_),
    .Y(_02352_));
 sky130_fd_sc_hd__a21oi_4 _08809_ (.A1(_02001_),
    .A2(_02183_),
    .B1(_02188_),
    .Y(_02353_));
 sky130_fd_sc_hd__and3_1 _08810_ (.A(_02351_),
    .B(_02352_),
    .C(_02353_),
    .X(_02354_));
 sky130_fd_sc_hd__a21oi_1 _08811_ (.A1(_02351_),
    .A2(_02352_),
    .B1(_02353_),
    .Y(_02355_));
 sky130_fd_sc_hd__or2_1 _08812_ (.A(_02354_),
    .B(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__a21oi_1 _08813_ (.A1(_02182_),
    .A2(_02187_),
    .B1(_02188_),
    .Y(_02357_));
 sky130_fd_sc_hd__or2_1 _08814_ (.A(_02356_),
    .B(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__xnor2_1 _08815_ (.A(_02356_),
    .B(_02357_),
    .Y(_02360_));
 sky130_fd_sc_hd__xor2_1 _08816_ (.A(_02346_),
    .B(_02360_),
    .X(_02361_));
 sky130_fd_sc_hd__o21a_1 _08817_ (.A1(_02178_),
    .A2(_02193_),
    .B1(_02192_),
    .X(_02362_));
 sky130_fd_sc_hd__and2b_1 _08818_ (.A_N(_02362_),
    .B(_02361_),
    .X(_02363_));
 sky130_fd_sc_hd__xnor2_1 _08819_ (.A(_02361_),
    .B(_02362_),
    .Y(_02364_));
 sky130_fd_sc_hd__xnor2_1 _08820_ (.A(_02334_),
    .B(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__a21oi_1 _08821_ (.A1(_02166_),
    .A2(_02198_),
    .B1(_02197_),
    .Y(_02366_));
 sky130_fd_sc_hd__nor2_1 _08822_ (.A(_02365_),
    .B(_02366_),
    .Y(_02367_));
 sky130_fd_sc_hd__xor2_1 _08823_ (.A(_02365_),
    .B(_02366_),
    .X(_02368_));
 sky130_fd_sc_hd__xor2_1 _08824_ (.A(_02311_),
    .B(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__a21oi_1 _08825_ (.A1(_02143_),
    .A2(_02202_),
    .B1(_02201_),
    .Y(_02371_));
 sky130_fd_sc_hd__and2b_1 _08826_ (.A_N(_02371_),
    .B(_02369_),
    .X(_02372_));
 sky130_fd_sc_hd__xnor2_1 _08827_ (.A(_02369_),
    .B(_02371_),
    .Y(_02373_));
 sky130_fd_sc_hd__xor2_1 _08828_ (.A(_02272_),
    .B(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__a21oi_1 _08829_ (.A1(_02103_),
    .A2(_02206_),
    .B1(_02205_),
    .Y(_02375_));
 sky130_fd_sc_hd__nand2b_1 _08830_ (.A_N(_02375_),
    .B(_02374_),
    .Y(_02376_));
 sky130_fd_sc_hd__xnor2_1 _08831_ (.A(_02374_),
    .B(_02375_),
    .Y(_02377_));
 sky130_fd_sc_hd__xnor2_1 _08832_ (.A(_02223_),
    .B(_02377_),
    .Y(_02378_));
 sky130_fd_sc_hd__a21oi_1 _08833_ (.A1(_02057_),
    .A2(_02210_),
    .B1(_02209_),
    .Y(_02379_));
 sky130_fd_sc_hd__or2_1 _08834_ (.A(_02378_),
    .B(_02379_),
    .X(_02380_));
 sky130_fd_sc_hd__xor2_1 _08835_ (.A(_02378_),
    .B(_02379_),
    .X(_02382_));
 sky130_fd_sc_hd__nand2_1 _08836_ (.A(_02222_),
    .B(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__xnor2_1 _08837_ (.A(_02222_),
    .B(_02382_),
    .Y(_02384_));
 sky130_fd_sc_hd__a21oi_2 _08838_ (.A1(_02056_),
    .A2(_02214_),
    .B1(_02213_),
    .Y(_02385_));
 sky130_fd_sc_hd__or2_1 _08839_ (.A(_02384_),
    .B(_02385_),
    .X(_02386_));
 sky130_fd_sc_hd__nand2_1 _08840_ (.A(_02384_),
    .B(_02385_),
    .Y(_02387_));
 sky130_fd_sc_hd__xnor2_1 _08841_ (.A(_02384_),
    .B(_02385_),
    .Y(_02388_));
 sky130_fd_sc_hd__o31a_1 _08842_ (.A1(_02040_),
    .A2(_02041_),
    .A3(_02219_),
    .B1(_02218_),
    .X(_02389_));
 sky130_fd_sc_hd__nor2_1 _08843_ (.A(_02042_),
    .B(_02220_),
    .Y(_02390_));
 sky130_fd_sc_hd__a21bo_1 _08844_ (.A1(_02053_),
    .A2(_02390_),
    .B1_N(_02389_),
    .X(_02391_));
 sky130_fd_sc_hd__xnor2_1 _08845_ (.A(_02388_),
    .B(_02391_),
    .Y(net92));
 sky130_fd_sc_hd__o21ai_1 _08846_ (.A1(_02070_),
    .A2(_02245_),
    .B1(_02244_),
    .Y(_02393_));
 sky130_fd_sc_hd__o21bai_1 _08847_ (.A1(_02225_),
    .A2(_02268_),
    .B1_N(_02270_),
    .Y(_02394_));
 sky130_fd_sc_hd__o21ba_1 _08848_ (.A1(_02246_),
    .A2(_02267_),
    .B1_N(_02266_),
    .X(_02395_));
 sky130_fd_sc_hd__a21boi_1 _08849_ (.A1(_02273_),
    .A2(_02310_),
    .B1_N(_02309_),
    .Y(_02396_));
 sky130_fd_sc_hd__and4_1 _08850_ (.A(net30),
    .B(net31),
    .C(net52),
    .D(net53),
    .X(_02397_));
 sky130_fd_sc_hd__a22oi_1 _08851_ (.A1(net31),
    .A2(net52),
    .B1(net53),
    .B2(net30),
    .Y(_02398_));
 sky130_fd_sc_hd__nor2_1 _08852_ (.A(_02397_),
    .B(_02398_),
    .Y(_02399_));
 sky130_fd_sc_hd__nand2_1 _08853_ (.A(net29),
    .B(net54),
    .Y(_02400_));
 sky130_fd_sc_hd__xnor2_1 _08854_ (.A(_02399_),
    .B(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__o21ba_1 _08855_ (.A1(_02228_),
    .A2(_02230_),
    .B1_N(_02226_),
    .X(_02403_));
 sky130_fd_sc_hd__nand2b_1 _08856_ (.A_N(_02403_),
    .B(_02401_),
    .Y(_02404_));
 sky130_fd_sc_hd__xnor2_1 _08857_ (.A(_02401_),
    .B(_02403_),
    .Y(_02405_));
 sky130_fd_sc_hd__and4b_1 _08858_ (.A_N(net27),
    .B(net56),
    .C(net57),
    .D(net28),
    .X(_02406_));
 sky130_fd_sc_hd__inv_2 _08859_ (.A(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__o2bb2a_1 _08860_ (.A1_N(net28),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net27),
    .X(_02408_));
 sky130_fd_sc_hd__nor2_1 _08861_ (.A(_02406_),
    .B(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__or2_1 _08862_ (.A(_02405_),
    .B(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__nand2_1 _08863_ (.A(_02405_),
    .B(_02409_),
    .Y(_02411_));
 sky130_fd_sc_hd__nand2_1 _08864_ (.A(_02410_),
    .B(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__nand2_1 _08865_ (.A(_02233_),
    .B(_02241_),
    .Y(_02414_));
 sky130_fd_sc_hd__nand2b_1 _08866_ (.A_N(_02412_),
    .B(_02414_),
    .Y(_02415_));
 sky130_fd_sc_hd__xor2_1 _08867_ (.A(_02412_),
    .B(_02414_),
    .X(_02416_));
 sky130_fd_sc_hd__xnor2_1 _08868_ (.A(_02236_),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__a21o_1 _08869_ (.A1(_02279_),
    .A2(_02288_),
    .B1(_02287_),
    .X(_02418_));
 sky130_fd_sc_hd__nand2_1 _08870_ (.A(_02251_),
    .B(_02254_),
    .Y(_02419_));
 sky130_fd_sc_hd__a31o_1 _08871_ (.A1(net3),
    .A2(net48),
    .A3(_02276_),
    .B1(_02275_),
    .X(_02420_));
 sky130_fd_sc_hd__nand4_2 _08872_ (.A(net2),
    .B(net3),
    .C(net49),
    .D(net50),
    .Y(_02421_));
 sky130_fd_sc_hd__a22o_1 _08873_ (.A1(net3),
    .A2(net49),
    .B1(net50),
    .B2(net2),
    .X(_02422_));
 sky130_fd_sc_hd__a22o_1 _08874_ (.A1(net32),
    .A2(net51),
    .B1(_02421_),
    .B2(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__nand4_2 _08875_ (.A(net32),
    .B(net51),
    .C(_02421_),
    .D(_02422_),
    .Y(_02425_));
 sky130_fd_sc_hd__nand3_2 _08876_ (.A(_02420_),
    .B(_02423_),
    .C(_02425_),
    .Y(_02426_));
 sky130_fd_sc_hd__a21o_1 _08877_ (.A1(_02423_),
    .A2(_02425_),
    .B1(_02420_),
    .X(_02427_));
 sky130_fd_sc_hd__nand3_2 _08878_ (.A(_02419_),
    .B(_02426_),
    .C(_02427_),
    .Y(_02428_));
 sky130_fd_sc_hd__a21o_1 _08879_ (.A1(_02426_),
    .A2(_02427_),
    .B1(_02419_),
    .X(_02429_));
 sky130_fd_sc_hd__and3_1 _08880_ (.A(_02418_),
    .B(_02428_),
    .C(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__a21oi_1 _08881_ (.A1(_02428_),
    .A2(_02429_),
    .B1(_02418_),
    .Y(_02431_));
 sky130_fd_sc_hd__a211oi_1 _08882_ (.A1(_02255_),
    .A2(_02257_),
    .B1(_02430_),
    .C1(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__o211a_1 _08883_ (.A1(_02430_),
    .A2(_02431_),
    .B1(_02255_),
    .C1(_02257_),
    .X(_02433_));
 sky130_fd_sc_hd__or2_1 _08884_ (.A(_02432_),
    .B(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__nor2_1 _08885_ (.A(_02259_),
    .B(_02262_),
    .Y(_02436_));
 sky130_fd_sc_hd__nor2_1 _08886_ (.A(_02434_),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__xnor2_1 _08887_ (.A(_02434_),
    .B(_02436_),
    .Y(_02438_));
 sky130_fd_sc_hd__xnor2_1 _08888_ (.A(_02417_),
    .B(_02438_),
    .Y(_02439_));
 sky130_fd_sc_hd__xor2_1 _08889_ (.A(_02396_),
    .B(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__and2b_1 _08890_ (.A_N(_02395_),
    .B(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__xnor2_1 _08891_ (.A(_02395_),
    .B(_02440_),
    .Y(_02442_));
 sky130_fd_sc_hd__nor2_1 _08892_ (.A(_02303_),
    .B(_02306_),
    .Y(_02443_));
 sky130_fd_sc_hd__and4_1 _08893_ (.A(net5),
    .B(net6),
    .C(net46),
    .D(net47),
    .X(_02444_));
 sky130_fd_sc_hd__a22o_1 _08894_ (.A1(net6),
    .A2(net46),
    .B1(net47),
    .B2(net5),
    .X(_02445_));
 sky130_fd_sc_hd__and2b_1 _08895_ (.A_N(_02444_),
    .B(_02445_),
    .X(_02447_));
 sky130_fd_sc_hd__nand2_1 _08896_ (.A(net4),
    .B(net48),
    .Y(_02448_));
 sky130_fd_sc_hd__xnor2_1 _08897_ (.A(_02447_),
    .B(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__nand2_1 _08898_ (.A(net7),
    .B(net45),
    .Y(_02450_));
 sky130_fd_sc_hd__and4_1 _08899_ (.A(net8),
    .B(net9),
    .C(net42),
    .D(net43),
    .X(_02451_));
 sky130_fd_sc_hd__a22oi_2 _08900_ (.A1(net9),
    .A2(net42),
    .B1(net43),
    .B2(net8),
    .Y(_02452_));
 sky130_fd_sc_hd__or3_1 _08901_ (.A(_02450_),
    .B(_02451_),
    .C(_02452_),
    .X(_02453_));
 sky130_fd_sc_hd__o21ai_1 _08902_ (.A1(_02451_),
    .A2(_02452_),
    .B1(_02450_),
    .Y(_02454_));
 sky130_fd_sc_hd__o21bai_1 _08903_ (.A1(_02280_),
    .A2(_02283_),
    .B1_N(_02281_),
    .Y(_02455_));
 sky130_fd_sc_hd__and3_1 _08904_ (.A(_02453_),
    .B(_02454_),
    .C(_02455_),
    .X(_02456_));
 sky130_fd_sc_hd__a21o_1 _08905_ (.A1(_02453_),
    .A2(_02454_),
    .B1(_02455_),
    .X(_02458_));
 sky130_fd_sc_hd__and2b_1 _08906_ (.A_N(_02456_),
    .B(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__xnor2_1 _08907_ (.A(_02449_),
    .B(_02459_),
    .Y(_02460_));
 sky130_fd_sc_hd__nand2_1 _08908_ (.A(_02294_),
    .B(_02297_),
    .Y(_02461_));
 sky130_fd_sc_hd__a31o_1 _08909_ (.A1(net38),
    .A2(net13),
    .A3(_02316_),
    .B1(_02314_),
    .X(_02462_));
 sky130_fd_sc_hd__nand4_1 _08910_ (.A(net39),
    .B(net40),
    .C(net11),
    .D(net13),
    .Y(_02463_));
 sky130_fd_sc_hd__a22o_1 _08911_ (.A1(net40),
    .A2(net11),
    .B1(net13),
    .B2(net39),
    .X(_02464_));
 sky130_fd_sc_hd__a22o_1 _08912_ (.A1(net41),
    .A2(net10),
    .B1(_02463_),
    .B2(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__nand4_1 _08913_ (.A(net41),
    .B(net10),
    .C(_02463_),
    .D(_02464_),
    .Y(_02466_));
 sky130_fd_sc_hd__nand3_1 _08914_ (.A(_02462_),
    .B(_02465_),
    .C(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__a21o_1 _08915_ (.A1(_02465_),
    .A2(_02466_),
    .B1(_02462_),
    .X(_02469_));
 sky130_fd_sc_hd__nand3_1 _08916_ (.A(_02461_),
    .B(_02467_),
    .C(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__a21o_1 _08917_ (.A1(_02467_),
    .A2(_02469_),
    .B1(_02461_),
    .X(_02471_));
 sky130_fd_sc_hd__a21bo_1 _08918_ (.A1(_02291_),
    .A2(_02299_),
    .B1_N(_02298_),
    .X(_02472_));
 sky130_fd_sc_hd__and3_1 _08919_ (.A(_02470_),
    .B(_02471_),
    .C(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__a21oi_1 _08920_ (.A1(_02470_),
    .A2(_02471_),
    .B1(_02472_),
    .Y(_02474_));
 sky130_fd_sc_hd__or3_1 _08921_ (.A(_02460_),
    .B(_02473_),
    .C(_02474_),
    .X(_02475_));
 sky130_fd_sc_hd__o21ai_1 _08922_ (.A1(_02473_),
    .A2(_02474_),
    .B1(_02460_),
    .Y(_02476_));
 sky130_fd_sc_hd__o211ai_1 _08923_ (.A1(_02330_),
    .A2(_02332_),
    .B1(_02475_),
    .C1(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__a211o_1 _08924_ (.A1(_02475_),
    .A2(_02476_),
    .B1(_02330_),
    .C1(_02332_),
    .X(_02478_));
 sky130_fd_sc_hd__nand2_1 _08925_ (.A(_02477_),
    .B(_02478_),
    .Y(_02480_));
 sky130_fd_sc_hd__xor2_1 _08926_ (.A(_02443_),
    .B(_02480_),
    .X(_02481_));
 sky130_fd_sc_hd__nand2_1 _08927_ (.A(_02325_),
    .B(_02328_),
    .Y(_02482_));
 sky130_fd_sc_hd__a21o_1 _08928_ (.A1(_02335_),
    .A2(_02344_),
    .B1(_02343_),
    .X(_02483_));
 sky130_fd_sc_hd__nand2_1 _08929_ (.A(net38),
    .B(net14),
    .Y(_02484_));
 sky130_fd_sc_hd__and4_1 _08930_ (.A(net36),
    .B(net37),
    .C(net15),
    .D(net16),
    .X(_02485_));
 sky130_fd_sc_hd__a22o_1 _08931_ (.A1(net37),
    .A2(net15),
    .B1(net16),
    .B2(net36),
    .X(_02486_));
 sky130_fd_sc_hd__and2b_1 _08932_ (.A_N(_02485_),
    .B(_02486_),
    .X(_02487_));
 sky130_fd_sc_hd__xnor2_1 _08933_ (.A(_02484_),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__nand2_1 _08934_ (.A(net35),
    .B(net17),
    .Y(_02489_));
 sky130_fd_sc_hd__and4_1 _08935_ (.A(net64),
    .B(net34),
    .C(net18),
    .D(net19),
    .X(_02491_));
 sky130_fd_sc_hd__a22oi_2 _08936_ (.A1(net34),
    .A2(net18),
    .B1(net19),
    .B2(net64),
    .Y(_02492_));
 sky130_fd_sc_hd__or3_1 _08937_ (.A(_02489_),
    .B(_02491_),
    .C(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__o21ai_1 _08938_ (.A1(_02491_),
    .A2(_02492_),
    .B1(_02489_),
    .Y(_02494_));
 sky130_fd_sc_hd__o21bai_1 _08939_ (.A1(_02319_),
    .A2(_02321_),
    .B1_N(_02320_),
    .Y(_02495_));
 sky130_fd_sc_hd__nand3_1 _08940_ (.A(_02493_),
    .B(_02494_),
    .C(_02495_),
    .Y(_02496_));
 sky130_fd_sc_hd__a21o_1 _08941_ (.A1(_02493_),
    .A2(_02494_),
    .B1(_02495_),
    .X(_02497_));
 sky130_fd_sc_hd__nand3_1 _08942_ (.A(_02488_),
    .B(_02496_),
    .C(_02497_),
    .Y(_02498_));
 sky130_fd_sc_hd__a21o_1 _08943_ (.A1(_02496_),
    .A2(_02497_),
    .B1(_02488_),
    .X(_02499_));
 sky130_fd_sc_hd__nand3_1 _08944_ (.A(_02483_),
    .B(_02498_),
    .C(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__a21o_1 _08945_ (.A1(_02498_),
    .A2(_02499_),
    .B1(_02483_),
    .X(_02502_));
 sky130_fd_sc_hd__and3_1 _08946_ (.A(_02482_),
    .B(_02500_),
    .C(_02502_),
    .X(_02503_));
 sky130_fd_sc_hd__a21oi_1 _08947_ (.A1(_02500_),
    .A2(_02502_),
    .B1(_02482_),
    .Y(_02504_));
 sky130_fd_sc_hd__nor2_1 _08948_ (.A(_02503_),
    .B(_02504_),
    .Y(_02505_));
 sky130_fd_sc_hd__nand2_1 _08949_ (.A(_02339_),
    .B(_02341_),
    .Y(_02506_));
 sky130_fd_sc_hd__o21bai_1 _08950_ (.A1(_02347_),
    .A2(_02350_),
    .B1_N(_02349_),
    .Y(_02507_));
 sky130_fd_sc_hd__a22o_1 _08951_ (.A1(net62),
    .A2(net21),
    .B1(net22),
    .B2(net61),
    .X(_02508_));
 sky130_fd_sc_hd__nand4_1 _08952_ (.A(net61),
    .B(net62),
    .C(net21),
    .D(net22),
    .Y(_02509_));
 sky130_fd_sc_hd__a22o_1 _08953_ (.A1(net63),
    .A2(net20),
    .B1(_02508_),
    .B2(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__nand4_1 _08954_ (.A(net63),
    .B(net20),
    .C(_02508_),
    .D(_02509_),
    .Y(_02511_));
 sky130_fd_sc_hd__nand3_1 _08955_ (.A(_02507_),
    .B(_02510_),
    .C(_02511_),
    .Y(_02513_));
 sky130_fd_sc_hd__a21o_1 _08956_ (.A1(_02510_),
    .A2(_02511_),
    .B1(_02507_),
    .X(_02514_));
 sky130_fd_sc_hd__and3_1 _08957_ (.A(_02506_),
    .B(_02513_),
    .C(_02514_),
    .X(_02515_));
 sky130_fd_sc_hd__a21oi_1 _08958_ (.A1(_02513_),
    .A2(_02514_),
    .B1(_02506_),
    .Y(_02516_));
 sky130_fd_sc_hd__and3_1 _08959_ (.A(net58),
    .B(net59),
    .C(net25),
    .X(_02517_));
 sky130_fd_sc_hd__nand3_1 _08960_ (.A(net58),
    .B(net59),
    .C(net25),
    .Y(_02518_));
 sky130_fd_sc_hd__o21a_1 _08961_ (.A1(net58),
    .A2(net59),
    .B1(net25),
    .X(_02519_));
 sky130_fd_sc_hd__a22o_1 _08962_ (.A1(net60),
    .A2(net24),
    .B1(_02518_),
    .B2(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__nand4_1 _08963_ (.A(net60),
    .B(net24),
    .C(_02518_),
    .D(_02519_),
    .Y(_02521_));
 sky130_fd_sc_hd__nand3_1 _08964_ (.A(_02353_),
    .B(_02520_),
    .C(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__a21o_1 _08965_ (.A1(_02520_),
    .A2(_02521_),
    .B1(_02353_),
    .X(_02524_));
 sky130_fd_sc_hd__a31o_1 _08966_ (.A1(_02351_),
    .A2(_02352_),
    .A3(_02353_),
    .B1(_02188_),
    .X(_02525_));
 sky130_fd_sc_hd__nand3_1 _08967_ (.A(_02522_),
    .B(_02524_),
    .C(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__a21o_1 _08968_ (.A1(_02522_),
    .A2(_02524_),
    .B1(_02525_),
    .X(_02527_));
 sky130_fd_sc_hd__or4bb_1 _08969_ (.A(_02515_),
    .B(_02516_),
    .C_N(_02526_),
    .D_N(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__a2bb2o_1 _08970_ (.A1_N(_02515_),
    .A2_N(_02516_),
    .B1(_02526_),
    .B2(_02527_),
    .X(_02529_));
 sky130_fd_sc_hd__nand2_1 _08971_ (.A(_02528_),
    .B(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__o21a_1 _08972_ (.A1(_02346_),
    .A2(_02360_),
    .B1(_02358_),
    .X(_02531_));
 sky130_fd_sc_hd__nor2_1 _08973_ (.A(_02530_),
    .B(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__xor2_1 _08974_ (.A(_02530_),
    .B(_02531_),
    .X(_02533_));
 sky130_fd_sc_hd__xnor2_1 _08975_ (.A(_02505_),
    .B(_02533_),
    .Y(_02535_));
 sky130_fd_sc_hd__a21oi_1 _08976_ (.A1(_02334_),
    .A2(_02364_),
    .B1(_02363_),
    .Y(_02536_));
 sky130_fd_sc_hd__nor2_1 _08977_ (.A(_02535_),
    .B(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__xor2_1 _08978_ (.A(_02535_),
    .B(_02536_),
    .X(_02538_));
 sky130_fd_sc_hd__xor2_1 _08979_ (.A(_02481_),
    .B(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__a21oi_1 _08980_ (.A1(_02311_),
    .A2(_02368_),
    .B1(_02367_),
    .Y(_02540_));
 sky130_fd_sc_hd__and2b_1 _08981_ (.A_N(_02540_),
    .B(_02539_),
    .X(_02541_));
 sky130_fd_sc_hd__xnor2_1 _08982_ (.A(_02539_),
    .B(_02540_),
    .Y(_02542_));
 sky130_fd_sc_hd__xor2_1 _08983_ (.A(_02442_),
    .B(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__a21oi_1 _08984_ (.A1(_02272_),
    .A2(_02373_),
    .B1(_02372_),
    .Y(_02544_));
 sky130_fd_sc_hd__nand2b_1 _08985_ (.A_N(_02544_),
    .B(_02543_),
    .Y(_02546_));
 sky130_fd_sc_hd__xnor2_1 _08986_ (.A(_02543_),
    .B(_02544_),
    .Y(_02547_));
 sky130_fd_sc_hd__xnor2_1 _08987_ (.A(_02394_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__a21boi_1 _08988_ (.A1(_02223_),
    .A2(_02377_),
    .B1_N(_02376_),
    .Y(_02549_));
 sky130_fd_sc_hd__nor2_1 _08989_ (.A(_02548_),
    .B(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__xor2_1 _08990_ (.A(_02548_),
    .B(_02549_),
    .X(_02551_));
 sky130_fd_sc_hd__xnor2_1 _08991_ (.A(_02393_),
    .B(_02551_),
    .Y(_02552_));
 sky130_fd_sc_hd__a21o_1 _08992_ (.A1(_02380_),
    .A2(_02383_),
    .B1(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__inv_2 _08993_ (.A(_02553_),
    .Y(_02554_));
 sky130_fd_sc_hd__and3_1 _08994_ (.A(_02380_),
    .B(_02383_),
    .C(_02552_),
    .X(_02555_));
 sky130_fd_sc_hd__nor2_1 _08995_ (.A(_02554_),
    .B(_02555_),
    .Y(_02557_));
 sky130_fd_sc_hd__a21boi_1 _08996_ (.A1(_02387_),
    .A2(_02391_),
    .B1_N(_02386_),
    .Y(_02558_));
 sky130_fd_sc_hd__xnor2_1 _08997_ (.A(_02557_),
    .B(_02558_),
    .Y(net93));
 sky130_fd_sc_hd__o21ai_1 _08998_ (.A1(_02236_),
    .A2(_02416_),
    .B1(_02415_),
    .Y(_02559_));
 sky130_fd_sc_hd__o21bai_1 _08999_ (.A1(_02396_),
    .A2(_02439_),
    .B1_N(_02441_),
    .Y(_02560_));
 sky130_fd_sc_hd__o21ba_1 _09000_ (.A1(_02417_),
    .A2(_02438_),
    .B1_N(_02437_),
    .X(_02561_));
 sky130_fd_sc_hd__o21ai_1 _09001_ (.A1(_02443_),
    .A2(_02480_),
    .B1(_02477_),
    .Y(_02562_));
 sky130_fd_sc_hd__and4_1 _09002_ (.A(net31),
    .B(net32),
    .C(net52),
    .D(net53),
    .X(_02563_));
 sky130_fd_sc_hd__a22o_1 _09003_ (.A1(net32),
    .A2(net52),
    .B1(net53),
    .B2(net31),
    .X(_02564_));
 sky130_fd_sc_hd__and2b_1 _09004_ (.A_N(_02563_),
    .B(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__nand2_1 _09005_ (.A(net30),
    .B(net54),
    .Y(_02567_));
 sky130_fd_sc_hd__xnor2_1 _09006_ (.A(_02565_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__o21ba_1 _09007_ (.A1(_02398_),
    .A2(_02400_),
    .B1_N(_02397_),
    .X(_02569_));
 sky130_fd_sc_hd__nand2b_1 _09008_ (.A_N(_02569_),
    .B(_02568_),
    .Y(_02570_));
 sky130_fd_sc_hd__xnor2_1 _09009_ (.A(_02568_),
    .B(_02569_),
    .Y(_02571_));
 sky130_fd_sc_hd__and4b_1 _09010_ (.A_N(net28),
    .B(net29),
    .C(net56),
    .D(net57),
    .X(_02572_));
 sky130_fd_sc_hd__inv_2 _09011_ (.A(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__o2bb2a_1 _09012_ (.A1_N(net29),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net28),
    .X(_02574_));
 sky130_fd_sc_hd__nor2_1 _09013_ (.A(_02572_),
    .B(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__or2_1 _09014_ (.A(_02571_),
    .B(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__nand2_1 _09015_ (.A(_02571_),
    .B(_02575_),
    .Y(_02578_));
 sky130_fd_sc_hd__nand2_1 _09016_ (.A(_02576_),
    .B(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__nand2_1 _09017_ (.A(_02404_),
    .B(_02411_),
    .Y(_02580_));
 sky130_fd_sc_hd__nand2b_1 _09018_ (.A_N(_02579_),
    .B(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__xor2_1 _09019_ (.A(_02579_),
    .B(_02580_),
    .X(_02582_));
 sky130_fd_sc_hd__xnor2_1 _09020_ (.A(_02407_),
    .B(_02582_),
    .Y(_02583_));
 sky130_fd_sc_hd__a21o_1 _09021_ (.A1(_02449_),
    .A2(_02458_),
    .B1(_02456_),
    .X(_02584_));
 sky130_fd_sc_hd__nand2_1 _09022_ (.A(_02421_),
    .B(_02425_),
    .Y(_02585_));
 sky130_fd_sc_hd__a31o_1 _09023_ (.A1(net4),
    .A2(net48),
    .A3(_02445_),
    .B1(_02444_),
    .X(_02586_));
 sky130_fd_sc_hd__nand4_2 _09024_ (.A(net3),
    .B(net4),
    .C(net49),
    .D(net50),
    .Y(_02587_));
 sky130_fd_sc_hd__a22o_1 _09025_ (.A1(net4),
    .A2(net49),
    .B1(net50),
    .B2(net3),
    .X(_02589_));
 sky130_fd_sc_hd__a22o_1 _09026_ (.A1(net2),
    .A2(net51),
    .B1(_02587_),
    .B2(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__nand4_2 _09027_ (.A(net2),
    .B(net51),
    .C(_02587_),
    .D(_02589_),
    .Y(_02591_));
 sky130_fd_sc_hd__nand3_2 _09028_ (.A(_02586_),
    .B(_02590_),
    .C(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__a21o_1 _09029_ (.A1(_02590_),
    .A2(_02591_),
    .B1(_02586_),
    .X(_02593_));
 sky130_fd_sc_hd__nand3_2 _09030_ (.A(_02585_),
    .B(_02592_),
    .C(_02593_),
    .Y(_02594_));
 sky130_fd_sc_hd__a21o_1 _09031_ (.A1(_02592_),
    .A2(_02593_),
    .B1(_02585_),
    .X(_02595_));
 sky130_fd_sc_hd__and3_1 _09032_ (.A(_02584_),
    .B(_02594_),
    .C(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__a21oi_1 _09033_ (.A1(_02594_),
    .A2(_02595_),
    .B1(_02584_),
    .Y(_02597_));
 sky130_fd_sc_hd__a211oi_1 _09034_ (.A1(_02426_),
    .A2(_02428_),
    .B1(_02596_),
    .C1(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__a211o_1 _09035_ (.A1(_02426_),
    .A2(_02428_),
    .B1(_02596_),
    .C1(_02597_),
    .X(_02600_));
 sky130_fd_sc_hd__o211ai_1 _09036_ (.A1(_02596_),
    .A2(_02597_),
    .B1(_02426_),
    .C1(_02428_),
    .Y(_02601_));
 sky130_fd_sc_hd__o211a_1 _09037_ (.A1(_02430_),
    .A2(_02432_),
    .B1(_02600_),
    .C1(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__a211oi_1 _09038_ (.A1(_02600_),
    .A2(_02601_),
    .B1(_02430_),
    .C1(_02432_),
    .Y(_02603_));
 sky130_fd_sc_hd__or2_1 _09039_ (.A(_02602_),
    .B(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__xnor2_1 _09040_ (.A(_02583_),
    .B(_02604_),
    .Y(_02605_));
 sky130_fd_sc_hd__and2b_1 _09041_ (.A_N(_02605_),
    .B(_02562_),
    .X(_02606_));
 sky130_fd_sc_hd__xnor2_1 _09042_ (.A(_02562_),
    .B(_02605_),
    .Y(_02607_));
 sky130_fd_sc_hd__and2b_1 _09043_ (.A_N(_02561_),
    .B(_02607_),
    .X(_02608_));
 sky130_fd_sc_hd__xnor2_1 _09044_ (.A(_02561_),
    .B(_02607_),
    .Y(_02609_));
 sky130_fd_sc_hd__and2b_1 _09045_ (.A_N(_02473_),
    .B(_02475_),
    .X(_02611_));
 sky130_fd_sc_hd__a21bo_1 _09046_ (.A1(_02482_),
    .A2(_02502_),
    .B1_N(_02500_),
    .X(_02612_));
 sky130_fd_sc_hd__and4_1 _09047_ (.A(net6),
    .B(net7),
    .C(net46),
    .D(net47),
    .X(_02613_));
 sky130_fd_sc_hd__a22o_1 _09048_ (.A1(net7),
    .A2(net46),
    .B1(net47),
    .B2(net6),
    .X(_02614_));
 sky130_fd_sc_hd__and2b_1 _09049_ (.A_N(_02613_),
    .B(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__nand2_1 _09050_ (.A(net5),
    .B(net48),
    .Y(_02616_));
 sky130_fd_sc_hd__xnor2_1 _09051_ (.A(_02615_),
    .B(_02616_),
    .Y(_02617_));
 sky130_fd_sc_hd__nand4_1 _09052_ (.A(net9),
    .B(net10),
    .C(net42),
    .D(net43),
    .Y(_02618_));
 sky130_fd_sc_hd__a22o_1 _09053_ (.A1(net10),
    .A2(net42),
    .B1(net43),
    .B2(net9),
    .X(_02619_));
 sky130_fd_sc_hd__and2_1 _09054_ (.A(net8),
    .B(net45),
    .X(_02620_));
 sky130_fd_sc_hd__a21o_1 _09055_ (.A1(_02618_),
    .A2(_02619_),
    .B1(_02620_),
    .X(_02622_));
 sky130_fd_sc_hd__nand3_1 _09056_ (.A(_02618_),
    .B(_02619_),
    .C(_02620_),
    .Y(_02623_));
 sky130_fd_sc_hd__o21bai_1 _09057_ (.A1(_02450_),
    .A2(_02452_),
    .B1_N(_02451_),
    .Y(_02624_));
 sky130_fd_sc_hd__and3_1 _09058_ (.A(_02622_),
    .B(_02623_),
    .C(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__a21o_1 _09059_ (.A1(_02622_),
    .A2(_02623_),
    .B1(_02624_),
    .X(_02626_));
 sky130_fd_sc_hd__and2b_1 _09060_ (.A_N(_02625_),
    .B(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__xnor2_1 _09061_ (.A(_02617_),
    .B(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__nand2_1 _09062_ (.A(_02463_),
    .B(_02466_),
    .Y(_02629_));
 sky130_fd_sc_hd__a31o_1 _09063_ (.A1(net38),
    .A2(net14),
    .A3(_02486_),
    .B1(_02485_),
    .X(_02630_));
 sky130_fd_sc_hd__nand4_1 _09064_ (.A(net39),
    .B(net40),
    .C(net13),
    .D(net14),
    .Y(_02631_));
 sky130_fd_sc_hd__a22o_1 _09065_ (.A1(net40),
    .A2(net13),
    .B1(net14),
    .B2(net39),
    .X(_02633_));
 sky130_fd_sc_hd__a22o_1 _09066_ (.A1(net41),
    .A2(net11),
    .B1(_02631_),
    .B2(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__nand4_1 _09067_ (.A(net41),
    .B(net11),
    .C(_02631_),
    .D(_02633_),
    .Y(_02635_));
 sky130_fd_sc_hd__nand3_1 _09068_ (.A(_02630_),
    .B(_02634_),
    .C(_02635_),
    .Y(_02636_));
 sky130_fd_sc_hd__a21o_1 _09069_ (.A1(_02634_),
    .A2(_02635_),
    .B1(_02630_),
    .X(_02637_));
 sky130_fd_sc_hd__nand3_1 _09070_ (.A(_02629_),
    .B(_02636_),
    .C(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__a21o_1 _09071_ (.A1(_02636_),
    .A2(_02637_),
    .B1(_02629_),
    .X(_02639_));
 sky130_fd_sc_hd__a21bo_1 _09072_ (.A1(_02461_),
    .A2(_02469_),
    .B1_N(_02467_),
    .X(_02640_));
 sky130_fd_sc_hd__and3_1 _09073_ (.A(_02638_),
    .B(_02639_),
    .C(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__inv_2 _09074_ (.A(_02641_),
    .Y(_02642_));
 sky130_fd_sc_hd__a21oi_1 _09075_ (.A1(_02638_),
    .A2(_02639_),
    .B1(_02640_),
    .Y(_02644_));
 sky130_fd_sc_hd__or3_1 _09076_ (.A(_02628_),
    .B(_02641_),
    .C(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__o21ai_1 _09077_ (.A1(_02641_),
    .A2(_02644_),
    .B1(_02628_),
    .Y(_02646_));
 sky130_fd_sc_hd__and3_1 _09078_ (.A(_02612_),
    .B(_02645_),
    .C(_02646_),
    .X(_02647_));
 sky130_fd_sc_hd__a21oi_1 _09079_ (.A1(_02645_),
    .A2(_02646_),
    .B1(_02612_),
    .Y(_02648_));
 sky130_fd_sc_hd__nor2_1 _09080_ (.A(_02647_),
    .B(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__xnor2_1 _09081_ (.A(_02611_),
    .B(_02649_),
    .Y(_02650_));
 sky130_fd_sc_hd__nand2_1 _09082_ (.A(_02496_),
    .B(_02498_),
    .Y(_02651_));
 sky130_fd_sc_hd__a21bo_1 _09083_ (.A1(_02506_),
    .A2(_02514_),
    .B1_N(_02513_),
    .X(_02652_));
 sky130_fd_sc_hd__and4_1 _09084_ (.A(net36),
    .B(net37),
    .C(net16),
    .D(net17),
    .X(_02653_));
 sky130_fd_sc_hd__a22o_1 _09085_ (.A1(net37),
    .A2(net16),
    .B1(net17),
    .B2(net36),
    .X(_02655_));
 sky130_fd_sc_hd__and2b_1 _09086_ (.A_N(_02653_),
    .B(_02655_),
    .X(_02656_));
 sky130_fd_sc_hd__nand2_1 _09087_ (.A(net38),
    .B(net15),
    .Y(_02657_));
 sky130_fd_sc_hd__xnor2_1 _09088_ (.A(_02656_),
    .B(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__nand4_1 _09089_ (.A(net64),
    .B(net34),
    .C(net19),
    .D(net20),
    .Y(_02659_));
 sky130_fd_sc_hd__a22o_1 _09090_ (.A1(net34),
    .A2(net19),
    .B1(net20),
    .B2(net64),
    .X(_02660_));
 sky130_fd_sc_hd__and2_1 _09091_ (.A(net35),
    .B(net18),
    .X(_02661_));
 sky130_fd_sc_hd__a21o_1 _09092_ (.A1(_02659_),
    .A2(_02660_),
    .B1(_02661_),
    .X(_02662_));
 sky130_fd_sc_hd__nand3_1 _09093_ (.A(_02659_),
    .B(_02660_),
    .C(_02661_),
    .Y(_02663_));
 sky130_fd_sc_hd__o21bai_1 _09094_ (.A1(_02489_),
    .A2(_02492_),
    .B1_N(_02491_),
    .Y(_02664_));
 sky130_fd_sc_hd__nand3_1 _09095_ (.A(_02662_),
    .B(_02663_),
    .C(_02664_),
    .Y(_02666_));
 sky130_fd_sc_hd__a21o_1 _09096_ (.A1(_02662_),
    .A2(_02663_),
    .B1(_02664_),
    .X(_02667_));
 sky130_fd_sc_hd__nand3_1 _09097_ (.A(_02658_),
    .B(_02666_),
    .C(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__a21o_1 _09098_ (.A1(_02666_),
    .A2(_02667_),
    .B1(_02658_),
    .X(_02669_));
 sky130_fd_sc_hd__nand3_2 _09099_ (.A(_02652_),
    .B(_02668_),
    .C(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__a21o_1 _09100_ (.A1(_02668_),
    .A2(_02669_),
    .B1(_02652_),
    .X(_02671_));
 sky130_fd_sc_hd__nand3_2 _09101_ (.A(_02651_),
    .B(_02670_),
    .C(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__a21o_1 _09102_ (.A1(_02670_),
    .A2(_02671_),
    .B1(_02651_),
    .X(_02673_));
 sky130_fd_sc_hd__nand2_1 _09103_ (.A(_02509_),
    .B(_02511_),
    .Y(_02674_));
 sky130_fd_sc_hd__a31o_1 _09104_ (.A1(net60),
    .A2(net24),
    .A3(_02519_),
    .B1(_02517_),
    .X(_02675_));
 sky130_fd_sc_hd__nand4_1 _09105_ (.A(net61),
    .B(net62),
    .C(net22),
    .D(net24),
    .Y(_02677_));
 sky130_fd_sc_hd__a22o_1 _09106_ (.A1(net62),
    .A2(net22),
    .B1(net24),
    .B2(net61),
    .X(_02678_));
 sky130_fd_sc_hd__a22o_1 _09107_ (.A1(net63),
    .A2(net21),
    .B1(_02677_),
    .B2(_02678_),
    .X(_02679_));
 sky130_fd_sc_hd__nand4_1 _09108_ (.A(net63),
    .B(net21),
    .C(_02677_),
    .D(_02678_),
    .Y(_02680_));
 sky130_fd_sc_hd__nand3_1 _09109_ (.A(_02675_),
    .B(_02679_),
    .C(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__a21o_1 _09110_ (.A1(_02679_),
    .A2(_02680_),
    .B1(_02675_),
    .X(_02682_));
 sky130_fd_sc_hd__nand3_1 _09111_ (.A(_02674_),
    .B(_02681_),
    .C(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__a21o_1 _09112_ (.A1(_02681_),
    .A2(_02682_),
    .B1(_02674_),
    .X(_02684_));
 sky130_fd_sc_hd__a22o_1 _09113_ (.A1(net60),
    .A2(net25),
    .B1(_02518_),
    .B2(_02519_),
    .X(_02685_));
 sky130_fd_sc_hd__nand4_1 _09114_ (.A(net60),
    .B(net25),
    .C(_02518_),
    .D(_02519_),
    .Y(_02686_));
 sky130_fd_sc_hd__a21o_1 _09115_ (.A1(_02685_),
    .A2(_02686_),
    .B1(_02353_),
    .X(_02688_));
 sky130_fd_sc_hd__nand3_1 _09116_ (.A(_02353_),
    .B(_02685_),
    .C(_02686_),
    .Y(_02689_));
 sky130_fd_sc_hd__a31o_1 _09117_ (.A1(_02353_),
    .A2(_02520_),
    .A3(_02521_),
    .B1(_02188_),
    .X(_02690_));
 sky130_fd_sc_hd__and3_1 _09118_ (.A(_02688_),
    .B(_02689_),
    .C(_02690_),
    .X(_02691_));
 sky130_fd_sc_hd__nand3_1 _09119_ (.A(_02688_),
    .B(_02689_),
    .C(_02690_),
    .Y(_02692_));
 sky130_fd_sc_hd__a21o_1 _09120_ (.A1(_02688_),
    .A2(_02689_),
    .B1(_02690_),
    .X(_02693_));
 sky130_fd_sc_hd__and4_1 _09121_ (.A(_02683_),
    .B(_02684_),
    .C(_02692_),
    .D(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__a22oi_2 _09122_ (.A1(_02683_),
    .A2(_02684_),
    .B1(_02692_),
    .B2(_02693_),
    .Y(_02695_));
 sky130_fd_sc_hd__a211o_1 _09123_ (.A1(_02526_),
    .A2(_02528_),
    .B1(_02694_),
    .C1(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__o211ai_2 _09124_ (.A1(_02694_),
    .A2(_02695_),
    .B1(_02526_),
    .C1(_02528_),
    .Y(_02697_));
 sky130_fd_sc_hd__nand4_1 _09125_ (.A(_02672_),
    .B(_02673_),
    .C(_02696_),
    .D(_02697_),
    .Y(_02699_));
 sky130_fd_sc_hd__a22o_1 _09126_ (.A1(_02672_),
    .A2(_02673_),
    .B1(_02696_),
    .B2(_02697_),
    .X(_02700_));
 sky130_fd_sc_hd__nand2_1 _09127_ (.A(_02699_),
    .B(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__a21oi_1 _09128_ (.A1(_02505_),
    .A2(_02533_),
    .B1(_02532_),
    .Y(_02702_));
 sky130_fd_sc_hd__nor2_1 _09129_ (.A(_02701_),
    .B(_02702_),
    .Y(_02703_));
 sky130_fd_sc_hd__xor2_1 _09130_ (.A(_02701_),
    .B(_02702_),
    .X(_02704_));
 sky130_fd_sc_hd__xor2_1 _09131_ (.A(_02650_),
    .B(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__a21oi_1 _09132_ (.A1(_02481_),
    .A2(_02538_),
    .B1(_02537_),
    .Y(_02706_));
 sky130_fd_sc_hd__and2b_1 _09133_ (.A_N(_02706_),
    .B(_02705_),
    .X(_02707_));
 sky130_fd_sc_hd__xnor2_1 _09134_ (.A(_02705_),
    .B(_02706_),
    .Y(_02708_));
 sky130_fd_sc_hd__xor2_1 _09135_ (.A(_02609_),
    .B(_02708_),
    .X(_02710_));
 sky130_fd_sc_hd__a21oi_1 _09136_ (.A1(_02442_),
    .A2(_02542_),
    .B1(_02541_),
    .Y(_02711_));
 sky130_fd_sc_hd__nand2b_1 _09137_ (.A_N(_02711_),
    .B(_02710_),
    .Y(_02712_));
 sky130_fd_sc_hd__xnor2_1 _09138_ (.A(_02710_),
    .B(_02711_),
    .Y(_02713_));
 sky130_fd_sc_hd__xnor2_1 _09139_ (.A(_02560_),
    .B(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__a21boi_1 _09140_ (.A1(_02394_),
    .A2(_02547_),
    .B1_N(_02546_),
    .Y(_02715_));
 sky130_fd_sc_hd__or2_1 _09141_ (.A(_02714_),
    .B(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__xor2_1 _09142_ (.A(_02714_),
    .B(_02715_),
    .X(_02717_));
 sky130_fd_sc_hd__nand2_1 _09143_ (.A(_02559_),
    .B(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__xnor2_1 _09144_ (.A(_02559_),
    .B(_02717_),
    .Y(_02719_));
 sky130_fd_sc_hd__a21oi_1 _09145_ (.A1(_02393_),
    .A2(_02551_),
    .B1(_02550_),
    .Y(_02721_));
 sky130_fd_sc_hd__or2_1 _09146_ (.A(_02719_),
    .B(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__nand2_1 _09147_ (.A(_02719_),
    .B(_02721_),
    .Y(_02723_));
 sky130_fd_sc_hd__nand2_1 _09148_ (.A(_02722_),
    .B(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__nor3_1 _09149_ (.A(_02388_),
    .B(_02554_),
    .C(_02555_),
    .Y(_02725_));
 sky130_fd_sc_hd__or3b_1 _09150_ (.A(_02555_),
    .B(_02388_),
    .C_N(_02553_),
    .X(_02726_));
 sky130_fd_sc_hd__o221ai_4 _09151_ (.A1(_02386_),
    .A2(_02555_),
    .B1(_02726_),
    .B2(_02389_),
    .C1(_02553_),
    .Y(_02727_));
 sky130_fd_sc_hd__a31o_1 _09152_ (.A1(_02053_),
    .A2(_02390_),
    .A3(_02725_),
    .B1(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__xnor2_1 _09153_ (.A(_02724_),
    .B(_02728_),
    .Y(net94));
 sky130_fd_sc_hd__o21ai_1 _09154_ (.A1(_02407_),
    .A2(_02582_),
    .B1(_02581_),
    .Y(_02729_));
 sky130_fd_sc_hd__or2_1 _09155_ (.A(_02606_),
    .B(_02608_),
    .X(_02731_));
 sky130_fd_sc_hd__o21ba_1 _09156_ (.A1(_02583_),
    .A2(_02604_),
    .B1_N(_02602_),
    .X(_02732_));
 sky130_fd_sc_hd__o21ba_1 _09157_ (.A1(_02611_),
    .A2(_02648_),
    .B1_N(_02647_),
    .X(_02733_));
 sky130_fd_sc_hd__and4_1 _09158_ (.A(net2),
    .B(net32),
    .C(net52),
    .D(net53),
    .X(_02734_));
 sky130_fd_sc_hd__a22o_1 _09159_ (.A1(net2),
    .A2(net52),
    .B1(net53),
    .B2(net32),
    .X(_02735_));
 sky130_fd_sc_hd__and2b_1 _09160_ (.A_N(_02734_),
    .B(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__nand2_1 _09161_ (.A(net31),
    .B(net54),
    .Y(_02737_));
 sky130_fd_sc_hd__xnor2_1 _09162_ (.A(_02736_),
    .B(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__a31o_1 _09163_ (.A1(net30),
    .A2(net54),
    .A3(_02564_),
    .B1(_02563_),
    .X(_02739_));
 sky130_fd_sc_hd__nand2_1 _09164_ (.A(_02738_),
    .B(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__xor2_1 _09165_ (.A(_02738_),
    .B(_02739_),
    .X(_02742_));
 sky130_fd_sc_hd__and4b_1 _09166_ (.A_N(net29),
    .B(net30),
    .C(net56),
    .D(net57),
    .X(_02743_));
 sky130_fd_sc_hd__o2bb2a_1 _09167_ (.A1_N(net30),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net29),
    .X(_02744_));
 sky130_fd_sc_hd__nor2_1 _09168_ (.A(_02743_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__xnor2_1 _09169_ (.A(_02742_),
    .B(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__nand3_1 _09170_ (.A(_02570_),
    .B(_02578_),
    .C(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__a21o_1 _09171_ (.A1(_02570_),
    .A2(_02578_),
    .B1(_02746_),
    .X(_02748_));
 sky130_fd_sc_hd__nand2_1 _09172_ (.A(_02747_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__xnor2_1 _09173_ (.A(_02573_),
    .B(_02749_),
    .Y(_02750_));
 sky130_fd_sc_hd__a21o_1 _09174_ (.A1(_02617_),
    .A2(_02626_),
    .B1(_02625_),
    .X(_02751_));
 sky130_fd_sc_hd__nand2_1 _09175_ (.A(_02587_),
    .B(_02591_),
    .Y(_02753_));
 sky130_fd_sc_hd__a31o_1 _09176_ (.A1(net5),
    .A2(net48),
    .A3(_02614_),
    .B1(_02613_),
    .X(_02754_));
 sky130_fd_sc_hd__nand4_2 _09177_ (.A(net4),
    .B(net5),
    .C(net49),
    .D(net50),
    .Y(_02755_));
 sky130_fd_sc_hd__a22o_1 _09178_ (.A1(net5),
    .A2(net49),
    .B1(net50),
    .B2(net4),
    .X(_02756_));
 sky130_fd_sc_hd__a22o_1 _09179_ (.A1(net3),
    .A2(net51),
    .B1(_02755_),
    .B2(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__nand4_2 _09180_ (.A(net3),
    .B(net51),
    .C(_02755_),
    .D(_02756_),
    .Y(_02758_));
 sky130_fd_sc_hd__nand3_2 _09181_ (.A(_02754_),
    .B(_02757_),
    .C(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__a21o_1 _09182_ (.A1(_02757_),
    .A2(_02758_),
    .B1(_02754_),
    .X(_02760_));
 sky130_fd_sc_hd__nand3_2 _09183_ (.A(_02753_),
    .B(_02759_),
    .C(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__a21o_1 _09184_ (.A1(_02759_),
    .A2(_02760_),
    .B1(_02753_),
    .X(_02762_));
 sky130_fd_sc_hd__and3_1 _09185_ (.A(_02751_),
    .B(_02761_),
    .C(_02762_),
    .X(_02764_));
 sky130_fd_sc_hd__a21oi_1 _09186_ (.A1(_02761_),
    .A2(_02762_),
    .B1(_02751_),
    .Y(_02765_));
 sky130_fd_sc_hd__a211oi_1 _09187_ (.A1(_02592_),
    .A2(_02594_),
    .B1(_02764_),
    .C1(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__a211o_1 _09188_ (.A1(_02592_),
    .A2(_02594_),
    .B1(_02764_),
    .C1(_02765_),
    .X(_02767_));
 sky130_fd_sc_hd__o211ai_1 _09189_ (.A1(_02764_),
    .A2(_02765_),
    .B1(_02592_),
    .C1(_02594_),
    .Y(_02768_));
 sky130_fd_sc_hd__o211a_1 _09190_ (.A1(_02596_),
    .A2(_02598_),
    .B1(_02767_),
    .C1(_02768_),
    .X(_02769_));
 sky130_fd_sc_hd__inv_2 _09191_ (.A(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__a211oi_1 _09192_ (.A1(_02767_),
    .A2(_02768_),
    .B1(_02596_),
    .C1(_02598_),
    .Y(_02771_));
 sky130_fd_sc_hd__nor2_1 _09193_ (.A(_02769_),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__or3_1 _09194_ (.A(_02750_),
    .B(_02769_),
    .C(_02771_),
    .X(_02773_));
 sky130_fd_sc_hd__xnor2_1 _09195_ (.A(_02750_),
    .B(_02772_),
    .Y(_02775_));
 sky130_fd_sc_hd__and2b_1 _09196_ (.A_N(_02733_),
    .B(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__xnor2_1 _09197_ (.A(_02733_),
    .B(_02775_),
    .Y(_02777_));
 sky130_fd_sc_hd__and2b_1 _09198_ (.A_N(_02732_),
    .B(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__xnor2_1 _09199_ (.A(_02732_),
    .B(_02777_),
    .Y(_02779_));
 sky130_fd_sc_hd__and4_1 _09200_ (.A(net7),
    .B(net8),
    .C(net46),
    .D(net47),
    .X(_02780_));
 sky130_fd_sc_hd__a22o_1 _09201_ (.A1(net8),
    .A2(net46),
    .B1(net47),
    .B2(net7),
    .X(_02781_));
 sky130_fd_sc_hd__and2b_1 _09202_ (.A_N(_02780_),
    .B(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__nand2_1 _09203_ (.A(net6),
    .B(net48),
    .Y(_02783_));
 sky130_fd_sc_hd__xnor2_2 _09204_ (.A(_02782_),
    .B(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__nand4_1 _09205_ (.A(net10),
    .B(net42),
    .C(net11),
    .D(net43),
    .Y(_02786_));
 sky130_fd_sc_hd__a22o_1 _09206_ (.A1(net42),
    .A2(net11),
    .B1(net43),
    .B2(net10),
    .X(_02787_));
 sky130_fd_sc_hd__and2_1 _09207_ (.A(net9),
    .B(net45),
    .X(_02788_));
 sky130_fd_sc_hd__a21o_1 _09208_ (.A1(_02786_),
    .A2(_02787_),
    .B1(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__nand3_1 _09209_ (.A(_02786_),
    .B(_02787_),
    .C(_02788_),
    .Y(_02790_));
 sky130_fd_sc_hd__a21bo_1 _09210_ (.A1(_02619_),
    .A2(_02620_),
    .B1_N(_02618_),
    .X(_02791_));
 sky130_fd_sc_hd__and3_1 _09211_ (.A(_02789_),
    .B(_02790_),
    .C(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__a21o_1 _09212_ (.A1(_02789_),
    .A2(_02790_),
    .B1(_02791_),
    .X(_02793_));
 sky130_fd_sc_hd__and2b_1 _09213_ (.A_N(_02792_),
    .B(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__xnor2_2 _09214_ (.A(_02784_),
    .B(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__nand2_1 _09215_ (.A(_02631_),
    .B(_02635_),
    .Y(_02797_));
 sky130_fd_sc_hd__a31o_1 _09216_ (.A1(net38),
    .A2(net15),
    .A3(_02655_),
    .B1(_02653_),
    .X(_02798_));
 sky130_fd_sc_hd__nand4_1 _09217_ (.A(net39),
    .B(net40),
    .C(net14),
    .D(net15),
    .Y(_02799_));
 sky130_fd_sc_hd__a22o_1 _09218_ (.A1(net40),
    .A2(net14),
    .B1(net15),
    .B2(net39),
    .X(_02800_));
 sky130_fd_sc_hd__a22o_1 _09219_ (.A1(net41),
    .A2(net13),
    .B1(_02799_),
    .B2(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__nand4_1 _09220_ (.A(net41),
    .B(net13),
    .C(_02799_),
    .D(_02800_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand3_1 _09221_ (.A(_02798_),
    .B(_02801_),
    .C(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__a21o_1 _09222_ (.A1(_02801_),
    .A2(_02802_),
    .B1(_02798_),
    .X(_02804_));
 sky130_fd_sc_hd__nand3_1 _09223_ (.A(_02797_),
    .B(_02803_),
    .C(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__a21o_1 _09224_ (.A1(_02803_),
    .A2(_02804_),
    .B1(_02797_),
    .X(_02806_));
 sky130_fd_sc_hd__a21bo_1 _09225_ (.A1(_02629_),
    .A2(_02637_),
    .B1_N(_02636_),
    .X(_02808_));
 sky130_fd_sc_hd__and3_1 _09226_ (.A(_02805_),
    .B(_02806_),
    .C(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__inv_2 _09227_ (.A(_02809_),
    .Y(_02810_));
 sky130_fd_sc_hd__a21oi_1 _09228_ (.A1(_02805_),
    .A2(_02806_),
    .B1(_02808_),
    .Y(_02811_));
 sky130_fd_sc_hd__nor3_1 _09229_ (.A(_02795_),
    .B(_02809_),
    .C(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__or3_1 _09230_ (.A(_02795_),
    .B(_02809_),
    .C(_02811_),
    .X(_02813_));
 sky130_fd_sc_hd__o21a_1 _09231_ (.A1(_02809_),
    .A2(_02811_),
    .B1(_02795_),
    .X(_02814_));
 sky130_fd_sc_hd__a211oi_2 _09232_ (.A1(_02670_),
    .A2(_02672_),
    .B1(_02812_),
    .C1(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__o211a_1 _09233_ (.A1(_02812_),
    .A2(_02814_),
    .B1(_02670_),
    .C1(_02672_),
    .X(_02816_));
 sky130_fd_sc_hd__a211oi_2 _09234_ (.A1(_02642_),
    .A2(_02645_),
    .B1(_02815_),
    .C1(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__o211a_1 _09235_ (.A1(_02815_),
    .A2(_02816_),
    .B1(_02642_),
    .C1(_02645_),
    .X(_02819_));
 sky130_fd_sc_hd__nand2_1 _09236_ (.A(_02666_),
    .B(_02668_),
    .Y(_02820_));
 sky130_fd_sc_hd__a21bo_1 _09237_ (.A1(_02674_),
    .A2(_02682_),
    .B1_N(_02681_),
    .X(_02821_));
 sky130_fd_sc_hd__and4_1 _09238_ (.A(net36),
    .B(net37),
    .C(net17),
    .D(net18),
    .X(_02822_));
 sky130_fd_sc_hd__a22o_1 _09239_ (.A1(net37),
    .A2(net17),
    .B1(net18),
    .B2(net36),
    .X(_02823_));
 sky130_fd_sc_hd__and2b_1 _09240_ (.A_N(_02822_),
    .B(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__nand2_1 _09241_ (.A(net38),
    .B(net16),
    .Y(_02825_));
 sky130_fd_sc_hd__xnor2_1 _09242_ (.A(_02824_),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__nand4_1 _09243_ (.A(net64),
    .B(net34),
    .C(net20),
    .D(net21),
    .Y(_02827_));
 sky130_fd_sc_hd__a22o_1 _09244_ (.A1(net34),
    .A2(net20),
    .B1(net21),
    .B2(net64),
    .X(_02828_));
 sky130_fd_sc_hd__and2_1 _09245_ (.A(net35),
    .B(net19),
    .X(_02830_));
 sky130_fd_sc_hd__a21o_1 _09246_ (.A1(_02827_),
    .A2(_02828_),
    .B1(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__nand3_1 _09247_ (.A(_02827_),
    .B(_02828_),
    .C(_02830_),
    .Y(_02832_));
 sky130_fd_sc_hd__a21bo_1 _09248_ (.A1(_02660_),
    .A2(_02661_),
    .B1_N(_02659_),
    .X(_02833_));
 sky130_fd_sc_hd__nand3_1 _09249_ (.A(_02831_),
    .B(_02832_),
    .C(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__a21o_1 _09250_ (.A1(_02831_),
    .A2(_02832_),
    .B1(_02833_),
    .X(_02835_));
 sky130_fd_sc_hd__nand3_1 _09251_ (.A(_02826_),
    .B(_02834_),
    .C(_02835_),
    .Y(_02836_));
 sky130_fd_sc_hd__a21o_1 _09252_ (.A1(_02834_),
    .A2(_02835_),
    .B1(_02826_),
    .X(_02837_));
 sky130_fd_sc_hd__nand3_2 _09253_ (.A(_02821_),
    .B(_02836_),
    .C(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__a21o_1 _09254_ (.A1(_02836_),
    .A2(_02837_),
    .B1(_02821_),
    .X(_02839_));
 sky130_fd_sc_hd__nand3_2 _09255_ (.A(_02820_),
    .B(_02838_),
    .C(_02839_),
    .Y(_02841_));
 sky130_fd_sc_hd__a21o_1 _09256_ (.A1(_02838_),
    .A2(_02839_),
    .B1(_02820_),
    .X(_02842_));
 sky130_fd_sc_hd__nand2_1 _09257_ (.A(_02677_),
    .B(_02680_),
    .Y(_02843_));
 sky130_fd_sc_hd__a31o_2 _09258_ (.A1(net60),
    .A2(net25),
    .A3(_02519_),
    .B1(_02517_),
    .X(_02844_));
 sky130_fd_sc_hd__nand4_1 _09259_ (.A(net61),
    .B(net62),
    .C(net24),
    .D(net25),
    .Y(_02845_));
 sky130_fd_sc_hd__a22o_1 _09260_ (.A1(net62),
    .A2(net24),
    .B1(net25),
    .B2(net61),
    .X(_02846_));
 sky130_fd_sc_hd__a22o_1 _09261_ (.A1(net63),
    .A2(net22),
    .B1(_02845_),
    .B2(_02846_),
    .X(_02847_));
 sky130_fd_sc_hd__nand4_1 _09262_ (.A(net63),
    .B(net22),
    .C(_02845_),
    .D(_02846_),
    .Y(_02848_));
 sky130_fd_sc_hd__nand3_1 _09263_ (.A(_02844_),
    .B(_02847_),
    .C(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__a21o_1 _09264_ (.A1(_02847_),
    .A2(_02848_),
    .B1(_02844_),
    .X(_02850_));
 sky130_fd_sc_hd__nand3_1 _09265_ (.A(_02843_),
    .B(_02849_),
    .C(_02850_),
    .Y(_02852_));
 sky130_fd_sc_hd__a21o_1 _09266_ (.A1(_02849_),
    .A2(_02850_),
    .B1(_02843_),
    .X(_02853_));
 sky130_fd_sc_hd__and3_1 _09267_ (.A(_02188_),
    .B(_02685_),
    .C(_02686_),
    .X(_02854_));
 sky130_fd_sc_hd__nor2_1 _09268_ (.A(_02188_),
    .B(_02688_),
    .Y(_02855_));
 sky130_fd_sc_hd__o21ba_2 _09269_ (.A1(_02188_),
    .A2(_02688_),
    .B1_N(_02854_),
    .X(_02856_));
 sky130_fd_sc_hd__nand3_1 _09270_ (.A(_02852_),
    .B(_02853_),
    .C(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__a21o_1 _09271_ (.A1(_02852_),
    .A2(_02853_),
    .B1(_02856_),
    .X(_02858_));
 sky130_fd_sc_hd__a31o_1 _09272_ (.A1(_02683_),
    .A2(_02684_),
    .A3(_02693_),
    .B1(_02691_),
    .X(_02859_));
 sky130_fd_sc_hd__nand3_2 _09273_ (.A(_02857_),
    .B(_02858_),
    .C(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__inv_2 _09274_ (.A(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__a21o_1 _09275_ (.A1(_02857_),
    .A2(_02858_),
    .B1(_02859_),
    .X(_02863_));
 sky130_fd_sc_hd__and4_1 _09276_ (.A(_02841_),
    .B(_02842_),
    .C(_02860_),
    .D(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__a22oi_2 _09277_ (.A1(_02841_),
    .A2(_02842_),
    .B1(_02860_),
    .B2(_02863_),
    .Y(_02865_));
 sky130_fd_sc_hd__a211o_1 _09278_ (.A1(_02696_),
    .A2(_02699_),
    .B1(_02864_),
    .C1(_02865_),
    .X(_02866_));
 sky130_fd_sc_hd__o211ai_1 _09279_ (.A1(_02864_),
    .A2(_02865_),
    .B1(_02696_),
    .C1(_02699_),
    .Y(_02867_));
 sky130_fd_sc_hd__or4bb_1 _09280_ (.A(_02817_),
    .B(_02819_),
    .C_N(_02866_),
    .D_N(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__a2bb2o_1 _09281_ (.A1_N(_02817_),
    .A2_N(_02819_),
    .B1(_02866_),
    .B2(_02867_),
    .X(_02869_));
 sky130_fd_sc_hd__nand2_1 _09282_ (.A(_02868_),
    .B(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__a21oi_1 _09283_ (.A1(_02650_),
    .A2(_02704_),
    .B1(_02703_),
    .Y(_02871_));
 sky130_fd_sc_hd__nor2_1 _09284_ (.A(_02870_),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__xor2_1 _09285_ (.A(_02870_),
    .B(_02871_),
    .X(_02874_));
 sky130_fd_sc_hd__xor2_1 _09286_ (.A(_02779_),
    .B(_02874_),
    .X(_02875_));
 sky130_fd_sc_hd__a21oi_1 _09287_ (.A1(_02609_),
    .A2(_02708_),
    .B1(_02707_),
    .Y(_02876_));
 sky130_fd_sc_hd__nand2b_1 _09288_ (.A_N(_02876_),
    .B(_02875_),
    .Y(_02877_));
 sky130_fd_sc_hd__xnor2_1 _09289_ (.A(_02875_),
    .B(_02876_),
    .Y(_02878_));
 sky130_fd_sc_hd__xnor2_1 _09290_ (.A(_02731_),
    .B(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__a21boi_1 _09291_ (.A1(_02560_),
    .A2(_02713_),
    .B1_N(_02712_),
    .Y(_02880_));
 sky130_fd_sc_hd__nor2_1 _09292_ (.A(_02879_),
    .B(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__xor2_1 _09293_ (.A(_02879_),
    .B(_02880_),
    .X(_02882_));
 sky130_fd_sc_hd__xnor2_1 _09294_ (.A(_02729_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__a21o_1 _09295_ (.A1(_02716_),
    .A2(_02718_),
    .B1(_02883_),
    .X(_02885_));
 sky130_fd_sc_hd__inv_2 _09296_ (.A(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__and3_1 _09297_ (.A(_02716_),
    .B(_02718_),
    .C(_02883_),
    .X(_02887_));
 sky130_fd_sc_hd__nor2_1 _09298_ (.A(_02886_),
    .B(_02887_),
    .Y(_02888_));
 sky130_fd_sc_hd__a21bo_1 _09299_ (.A1(_02723_),
    .A2(_02728_),
    .B1_N(_02722_),
    .X(_02889_));
 sky130_fd_sc_hd__xor2_1 _09300_ (.A(_02888_),
    .B(_02889_),
    .X(net95));
 sky130_fd_sc_hd__o21ai_1 _09301_ (.A1(_02573_),
    .A2(_02749_),
    .B1(_02748_),
    .Y(_02890_));
 sky130_fd_sc_hd__or2_1 _09302_ (.A(_02776_),
    .B(_02778_),
    .X(_02891_));
 sky130_fd_sc_hd__and4_1 _09303_ (.A(net2),
    .B(net3),
    .C(net52),
    .D(net53),
    .X(_02892_));
 sky130_fd_sc_hd__a22o_1 _09304_ (.A1(net3),
    .A2(net52),
    .B1(net53),
    .B2(net2),
    .X(_02893_));
 sky130_fd_sc_hd__and2b_1 _09305_ (.A_N(_02892_),
    .B(_02893_),
    .X(_02895_));
 sky130_fd_sc_hd__nand2_1 _09306_ (.A(net32),
    .B(net54),
    .Y(_02896_));
 sky130_fd_sc_hd__xnor2_1 _09307_ (.A(_02895_),
    .B(_02896_),
    .Y(_02897_));
 sky130_fd_sc_hd__a31o_1 _09308_ (.A1(net31),
    .A2(net54),
    .A3(_02735_),
    .B1(_02734_),
    .X(_02898_));
 sky130_fd_sc_hd__nand2_1 _09309_ (.A(_02897_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__xor2_1 _09310_ (.A(_02897_),
    .B(_02898_),
    .X(_02900_));
 sky130_fd_sc_hd__and4b_1 _09311_ (.A_N(net30),
    .B(net31),
    .C(net56),
    .D(net57),
    .X(_02901_));
 sky130_fd_sc_hd__o2bb2a_1 _09312_ (.A1_N(net31),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net30),
    .X(_02902_));
 sky130_fd_sc_hd__nor2_1 _09313_ (.A(_02901_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__xnor2_1 _09314_ (.A(_02900_),
    .B(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__a21bo_1 _09315_ (.A1(_02742_),
    .A2(_02745_),
    .B1_N(_02740_),
    .X(_02906_));
 sky130_fd_sc_hd__and2b_1 _09316_ (.A_N(_02904_),
    .B(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__xor2_1 _09317_ (.A(_02904_),
    .B(_02906_),
    .X(_02908_));
 sky130_fd_sc_hd__inv_2 _09318_ (.A(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__xor2_1 _09319_ (.A(_02743_),
    .B(_02908_),
    .X(_02910_));
 sky130_fd_sc_hd__a21o_1 _09320_ (.A1(_02784_),
    .A2(_02793_),
    .B1(_02792_),
    .X(_02911_));
 sky130_fd_sc_hd__nand2_1 _09321_ (.A(_02755_),
    .B(_02758_),
    .Y(_02912_));
 sky130_fd_sc_hd__a31o_1 _09322_ (.A1(net6),
    .A2(net48),
    .A3(_02781_),
    .B1(_02780_),
    .X(_02913_));
 sky130_fd_sc_hd__nand4_2 _09323_ (.A(net5),
    .B(net6),
    .C(net49),
    .D(net50),
    .Y(_02914_));
 sky130_fd_sc_hd__a22o_1 _09324_ (.A1(net6),
    .A2(net49),
    .B1(net50),
    .B2(net5),
    .X(_02915_));
 sky130_fd_sc_hd__a22o_1 _09325_ (.A1(net4),
    .A2(net51),
    .B1(_02914_),
    .B2(_02915_),
    .X(_02917_));
 sky130_fd_sc_hd__nand4_2 _09326_ (.A(net4),
    .B(net51),
    .C(_02914_),
    .D(_02915_),
    .Y(_02918_));
 sky130_fd_sc_hd__nand3_2 _09327_ (.A(_02913_),
    .B(_02917_),
    .C(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__a21o_1 _09328_ (.A1(_02917_),
    .A2(_02918_),
    .B1(_02913_),
    .X(_02920_));
 sky130_fd_sc_hd__nand3_2 _09329_ (.A(_02912_),
    .B(_02919_),
    .C(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__a21o_1 _09330_ (.A1(_02919_),
    .A2(_02920_),
    .B1(_02912_),
    .X(_02922_));
 sky130_fd_sc_hd__and3_1 _09331_ (.A(_02911_),
    .B(_02921_),
    .C(_02922_),
    .X(_02923_));
 sky130_fd_sc_hd__a21oi_1 _09332_ (.A1(_02921_),
    .A2(_02922_),
    .B1(_02911_),
    .Y(_02924_));
 sky130_fd_sc_hd__a211oi_1 _09333_ (.A1(_02759_),
    .A2(_02761_),
    .B1(_02923_),
    .C1(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__a211o_1 _09334_ (.A1(_02759_),
    .A2(_02761_),
    .B1(_02923_),
    .C1(_02924_),
    .X(_02926_));
 sky130_fd_sc_hd__o211ai_1 _09335_ (.A1(_02923_),
    .A2(_02924_),
    .B1(_02759_),
    .C1(_02761_),
    .Y(_02928_));
 sky130_fd_sc_hd__o211a_1 _09336_ (.A1(_02764_),
    .A2(_02766_),
    .B1(_02926_),
    .C1(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__inv_2 _09337_ (.A(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__a211oi_1 _09338_ (.A1(_02926_),
    .A2(_02928_),
    .B1(_02764_),
    .C1(_02766_),
    .Y(_02931_));
 sky130_fd_sc_hd__or3_2 _09339_ (.A(_02910_),
    .B(_02929_),
    .C(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__o21ai_1 _09340_ (.A1(_02929_),
    .A2(_02931_),
    .B1(_02910_),
    .Y(_02933_));
 sky130_fd_sc_hd__o211a_1 _09341_ (.A1(_02815_),
    .A2(_02817_),
    .B1(_02932_),
    .C1(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__a211oi_1 _09342_ (.A1(_02932_),
    .A2(_02933_),
    .B1(_02815_),
    .C1(_02817_),
    .Y(_02935_));
 sky130_fd_sc_hd__a211oi_1 _09343_ (.A1(_02770_),
    .A2(_02773_),
    .B1(_02934_),
    .C1(_02935_),
    .Y(_02936_));
 sky130_fd_sc_hd__o211a_1 _09344_ (.A1(_02934_),
    .A2(_02935_),
    .B1(_02770_),
    .C1(_02773_),
    .X(_02937_));
 sky130_fd_sc_hd__and4_1 _09345_ (.A(net8),
    .B(net9),
    .C(net46),
    .D(net47),
    .X(_02939_));
 sky130_fd_sc_hd__a22o_1 _09346_ (.A1(net9),
    .A2(net46),
    .B1(net47),
    .B2(net8),
    .X(_02940_));
 sky130_fd_sc_hd__and2b_1 _09347_ (.A_N(_02939_),
    .B(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__nand2_1 _09348_ (.A(net7),
    .B(net48),
    .Y(_02942_));
 sky130_fd_sc_hd__xnor2_2 _09349_ (.A(_02941_),
    .B(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__nand4_1 _09350_ (.A(net42),
    .B(net11),
    .C(net43),
    .D(net13),
    .Y(_02944_));
 sky130_fd_sc_hd__a22o_1 _09351_ (.A1(net11),
    .A2(net43),
    .B1(net13),
    .B2(net42),
    .X(_02945_));
 sky130_fd_sc_hd__and2_1 _09352_ (.A(net10),
    .B(net45),
    .X(_02946_));
 sky130_fd_sc_hd__a21o_1 _09353_ (.A1(_02944_),
    .A2(_02945_),
    .B1(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__nand3_1 _09354_ (.A(_02944_),
    .B(_02945_),
    .C(_02946_),
    .Y(_02948_));
 sky130_fd_sc_hd__a21bo_1 _09355_ (.A1(_02787_),
    .A2(_02788_),
    .B1_N(_02786_),
    .X(_02950_));
 sky130_fd_sc_hd__and3_1 _09356_ (.A(_02947_),
    .B(_02948_),
    .C(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__a21o_1 _09357_ (.A1(_02947_),
    .A2(_02948_),
    .B1(_02950_),
    .X(_02952_));
 sky130_fd_sc_hd__and2b_1 _09358_ (.A_N(_02951_),
    .B(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__xnor2_2 _09359_ (.A(_02943_),
    .B(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__nand2_1 _09360_ (.A(_02799_),
    .B(_02802_),
    .Y(_02955_));
 sky130_fd_sc_hd__a31o_1 _09361_ (.A1(net38),
    .A2(net16),
    .A3(_02823_),
    .B1(_02822_),
    .X(_02956_));
 sky130_fd_sc_hd__nand4_1 _09362_ (.A(net39),
    .B(net40),
    .C(net15),
    .D(net16),
    .Y(_02957_));
 sky130_fd_sc_hd__a22o_1 _09363_ (.A1(net40),
    .A2(net15),
    .B1(net16),
    .B2(net39),
    .X(_02958_));
 sky130_fd_sc_hd__a22o_1 _09364_ (.A1(net41),
    .A2(net14),
    .B1(_02957_),
    .B2(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__nand4_1 _09365_ (.A(net41),
    .B(net14),
    .C(_02957_),
    .D(_02958_),
    .Y(_02961_));
 sky130_fd_sc_hd__nand3_1 _09366_ (.A(_02956_),
    .B(_02959_),
    .C(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__a21o_1 _09367_ (.A1(_02959_),
    .A2(_02961_),
    .B1(_02956_),
    .X(_02963_));
 sky130_fd_sc_hd__nand3_1 _09368_ (.A(_02955_),
    .B(_02962_),
    .C(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hd__a21o_1 _09369_ (.A1(_02962_),
    .A2(_02963_),
    .B1(_02955_),
    .X(_02965_));
 sky130_fd_sc_hd__a21bo_1 _09370_ (.A1(_02797_),
    .A2(_02804_),
    .B1_N(_02803_),
    .X(_02966_));
 sky130_fd_sc_hd__and3_1 _09371_ (.A(_02964_),
    .B(_02965_),
    .C(_02966_),
    .X(_02967_));
 sky130_fd_sc_hd__inv_2 _09372_ (.A(_02967_),
    .Y(_02968_));
 sky130_fd_sc_hd__a21oi_1 _09373_ (.A1(_02964_),
    .A2(_02965_),
    .B1(_02966_),
    .Y(_02969_));
 sky130_fd_sc_hd__nor3_1 _09374_ (.A(_02954_),
    .B(_02967_),
    .C(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__or3_1 _09375_ (.A(_02954_),
    .B(_02967_),
    .C(_02969_),
    .X(_02972_));
 sky130_fd_sc_hd__o21a_1 _09376_ (.A1(_02967_),
    .A2(_02969_),
    .B1(_02954_),
    .X(_02973_));
 sky130_fd_sc_hd__a211oi_4 _09377_ (.A1(_02838_),
    .A2(_02841_),
    .B1(_02970_),
    .C1(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__o211a_1 _09378_ (.A1(_02970_),
    .A2(_02973_),
    .B1(_02838_),
    .C1(_02841_),
    .X(_02975_));
 sky130_fd_sc_hd__a211oi_2 _09379_ (.A1(_02810_),
    .A2(_02813_),
    .B1(_02974_),
    .C1(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__o211a_1 _09380_ (.A1(_02974_),
    .A2(_02975_),
    .B1(_02810_),
    .C1(_02813_),
    .X(_02977_));
 sky130_fd_sc_hd__nand2_1 _09381_ (.A(_02834_),
    .B(_02836_),
    .Y(_02978_));
 sky130_fd_sc_hd__a21bo_1 _09382_ (.A1(_02843_),
    .A2(_02850_),
    .B1_N(_02849_),
    .X(_02979_));
 sky130_fd_sc_hd__and4_1 _09383_ (.A(net36),
    .B(net37),
    .C(net18),
    .D(net19),
    .X(_02980_));
 sky130_fd_sc_hd__a22o_1 _09384_ (.A1(net37),
    .A2(net18),
    .B1(net19),
    .B2(net36),
    .X(_02981_));
 sky130_fd_sc_hd__and2b_1 _09385_ (.A_N(_02980_),
    .B(_02981_),
    .X(_02983_));
 sky130_fd_sc_hd__nand2_1 _09386_ (.A(net38),
    .B(net17),
    .Y(_02984_));
 sky130_fd_sc_hd__xnor2_1 _09387_ (.A(_02983_),
    .B(_02984_),
    .Y(_02985_));
 sky130_fd_sc_hd__nand4_1 _09388_ (.A(net64),
    .B(net34),
    .C(net21),
    .D(net22),
    .Y(_02986_));
 sky130_fd_sc_hd__a22o_1 _09389_ (.A1(net34),
    .A2(net21),
    .B1(net22),
    .B2(net64),
    .X(_02987_));
 sky130_fd_sc_hd__and2_1 _09390_ (.A(net35),
    .B(net20),
    .X(_02988_));
 sky130_fd_sc_hd__a21o_1 _09391_ (.A1(_02986_),
    .A2(_02987_),
    .B1(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__nand3_1 _09392_ (.A(_02986_),
    .B(_02987_),
    .C(_02988_),
    .Y(_02990_));
 sky130_fd_sc_hd__a21bo_1 _09393_ (.A1(_02828_),
    .A2(_02830_),
    .B1_N(_02827_),
    .X(_02991_));
 sky130_fd_sc_hd__nand3_1 _09394_ (.A(_02989_),
    .B(_02990_),
    .C(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__a21o_1 _09395_ (.A1(_02989_),
    .A2(_02990_),
    .B1(_02991_),
    .X(_02994_));
 sky130_fd_sc_hd__nand3_1 _09396_ (.A(_02985_),
    .B(_02992_),
    .C(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__a21o_1 _09397_ (.A1(_02992_),
    .A2(_02994_),
    .B1(_02985_),
    .X(_02996_));
 sky130_fd_sc_hd__nand3_2 _09398_ (.A(_02979_),
    .B(_02995_),
    .C(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__a21o_1 _09399_ (.A1(_02995_),
    .A2(_02996_),
    .B1(_02979_),
    .X(_02998_));
 sky130_fd_sc_hd__nand3_2 _09400_ (.A(_02978_),
    .B(_02997_),
    .C(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__a21o_1 _09401_ (.A1(_02997_),
    .A2(_02998_),
    .B1(_02978_),
    .X(_03000_));
 sky130_fd_sc_hd__nand2_1 _09402_ (.A(_02845_),
    .B(_02848_),
    .Y(_03001_));
 sky130_fd_sc_hd__nand3_2 _09403_ (.A(net61),
    .B(net62),
    .C(net25),
    .Y(_03002_));
 sky130_fd_sc_hd__o21a_1 _09404_ (.A1(net61),
    .A2(net62),
    .B1(net25),
    .X(_03003_));
 sky130_fd_sc_hd__a22o_1 _09405_ (.A1(net63),
    .A2(net24),
    .B1(_03002_),
    .B2(_03003_),
    .X(_03005_));
 sky130_fd_sc_hd__nand4_1 _09406_ (.A(net63),
    .B(net24),
    .C(_03002_),
    .D(_03003_),
    .Y(_03006_));
 sky130_fd_sc_hd__nand3_1 _09407_ (.A(_02844_),
    .B(_03005_),
    .C(_03006_),
    .Y(_03007_));
 sky130_fd_sc_hd__a21o_1 _09408_ (.A1(_03005_),
    .A2(_03006_),
    .B1(_02844_),
    .X(_03008_));
 sky130_fd_sc_hd__nand3_1 _09409_ (.A(_03001_),
    .B(_03007_),
    .C(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__a21o_1 _09410_ (.A1(_03007_),
    .A2(_03008_),
    .B1(_03001_),
    .X(_03010_));
 sky130_fd_sc_hd__nand3_1 _09411_ (.A(_02856_),
    .B(_03009_),
    .C(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__a21o_1 _09412_ (.A1(_03009_),
    .A2(_03010_),
    .B1(_02856_),
    .X(_03012_));
 sky130_fd_sc_hd__a31o_1 _09413_ (.A1(_02852_),
    .A2(_02853_),
    .A3(_02856_),
    .B1(_02854_),
    .X(_03013_));
 sky130_fd_sc_hd__nand3_2 _09414_ (.A(_03011_),
    .B(_03012_),
    .C(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__inv_2 _09415_ (.A(_03014_),
    .Y(_03016_));
 sky130_fd_sc_hd__a21o_1 _09416_ (.A1(_03011_),
    .A2(_03012_),
    .B1(_03013_),
    .X(_03017_));
 sky130_fd_sc_hd__and4_1 _09417_ (.A(_02999_),
    .B(_03000_),
    .C(_03014_),
    .D(_03017_),
    .X(_03018_));
 sky130_fd_sc_hd__nand4_1 _09418_ (.A(_02999_),
    .B(_03000_),
    .C(_03014_),
    .D(_03017_),
    .Y(_03019_));
 sky130_fd_sc_hd__a22o_1 _09419_ (.A1(_02999_),
    .A2(_03000_),
    .B1(_03014_),
    .B2(_03017_),
    .X(_03020_));
 sky130_fd_sc_hd__o211a_1 _09420_ (.A1(_02861_),
    .A2(_02864_),
    .B1(_03019_),
    .C1(_03020_),
    .X(_03021_));
 sky130_fd_sc_hd__a211oi_2 _09421_ (.A1(_03019_),
    .A2(_03020_),
    .B1(_02861_),
    .C1(_02864_),
    .Y(_03022_));
 sky130_fd_sc_hd__nor4_2 _09422_ (.A(_02976_),
    .B(_02977_),
    .C(_03021_),
    .D(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__o22a_1 _09423_ (.A1(_02976_),
    .A2(_02977_),
    .B1(_03021_),
    .B2(_03022_),
    .X(_03024_));
 sky130_fd_sc_hd__a211oi_2 _09424_ (.A1(_02866_),
    .A2(_02868_),
    .B1(_03023_),
    .C1(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__o211a_1 _09425_ (.A1(_03023_),
    .A2(_03024_),
    .B1(_02866_),
    .C1(_02868_),
    .X(_03027_));
 sky130_fd_sc_hd__nor4_1 _09426_ (.A(_02936_),
    .B(_02937_),
    .C(_03025_),
    .D(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__o22a_1 _09427_ (.A1(_02936_),
    .A2(_02937_),
    .B1(_03025_),
    .B2(_03027_),
    .X(_03029_));
 sky130_fd_sc_hd__or2_1 _09428_ (.A(_03028_),
    .B(_03029_),
    .X(_03030_));
 sky130_fd_sc_hd__a21oi_1 _09429_ (.A1(_02779_),
    .A2(_02874_),
    .B1(_02872_),
    .Y(_03031_));
 sky130_fd_sc_hd__nor2_1 _09430_ (.A(_03030_),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__xor2_1 _09431_ (.A(_03030_),
    .B(_03031_),
    .X(_03033_));
 sky130_fd_sc_hd__xnor2_1 _09432_ (.A(_02891_),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__a21boi_1 _09433_ (.A1(_02731_),
    .A2(_02878_),
    .B1_N(_02877_),
    .Y(_03035_));
 sky130_fd_sc_hd__nor2_1 _09434_ (.A(_03034_),
    .B(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__xor2_1 _09435_ (.A(_03034_),
    .B(_03035_),
    .X(_03038_));
 sky130_fd_sc_hd__xnor2_1 _09436_ (.A(_02890_),
    .B(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__a21oi_1 _09437_ (.A1(_02729_),
    .A2(_02882_),
    .B1(_02881_),
    .Y(_03040_));
 sky130_fd_sc_hd__or2_1 _09438_ (.A(_03039_),
    .B(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__nand2_1 _09439_ (.A(_03039_),
    .B(_03040_),
    .Y(_03042_));
 sky130_fd_sc_hd__xnor2_1 _09440_ (.A(_03039_),
    .B(_03040_),
    .Y(_03043_));
 sky130_fd_sc_hd__a21oi_1 _09441_ (.A1(_02722_),
    .A2(_02885_),
    .B1(_02887_),
    .Y(_03044_));
 sky130_fd_sc_hd__nor3_2 _09442_ (.A(_02724_),
    .B(_02886_),
    .C(_02887_),
    .Y(_03045_));
 sky130_fd_sc_hd__a21o_1 _09443_ (.A1(_02728_),
    .A2(_03045_),
    .B1(_03044_),
    .X(_03046_));
 sky130_fd_sc_hd__xnor2_1 _09444_ (.A(_03043_),
    .B(_03046_),
    .Y(net96));
 sky130_fd_sc_hd__a21oi_1 _09445_ (.A1(_02890_),
    .A2(_03038_),
    .B1(_03036_),
    .Y(_03048_));
 sky130_fd_sc_hd__a21o_1 _09446_ (.A1(_02743_),
    .A2(_02909_),
    .B1(_02907_),
    .X(_03049_));
 sky130_fd_sc_hd__nor2_1 _09447_ (.A(_02934_),
    .B(_02936_),
    .Y(_03050_));
 sky130_fd_sc_hd__and4_1 _09448_ (.A(net3),
    .B(net4),
    .C(net52),
    .D(net53),
    .X(_03051_));
 sky130_fd_sc_hd__a22o_1 _09449_ (.A1(net4),
    .A2(net52),
    .B1(net53),
    .B2(net3),
    .X(_03052_));
 sky130_fd_sc_hd__and2b_1 _09450_ (.A_N(_03051_),
    .B(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__nand2_1 _09451_ (.A(net2),
    .B(net54),
    .Y(_03054_));
 sky130_fd_sc_hd__xnor2_1 _09452_ (.A(_03053_),
    .B(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__a31o_1 _09453_ (.A1(net32),
    .A2(net54),
    .A3(_02893_),
    .B1(_02892_),
    .X(_03056_));
 sky130_fd_sc_hd__nand2_1 _09454_ (.A(_03055_),
    .B(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__xor2_1 _09455_ (.A(_03055_),
    .B(_03056_),
    .X(_03059_));
 sky130_fd_sc_hd__and4b_1 _09456_ (.A_N(net31),
    .B(net32),
    .C(net56),
    .D(net57),
    .X(_03060_));
 sky130_fd_sc_hd__o2bb2a_1 _09457_ (.A1_N(net32),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net31),
    .X(_03061_));
 sky130_fd_sc_hd__nor2_1 _09458_ (.A(_03060_),
    .B(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__xnor2_1 _09459_ (.A(_03059_),
    .B(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__a21bo_1 _09460_ (.A1(_02900_),
    .A2(_02903_),
    .B1_N(_02899_),
    .X(_03064_));
 sky130_fd_sc_hd__and2b_1 _09461_ (.A_N(_03063_),
    .B(_03064_),
    .X(_03065_));
 sky130_fd_sc_hd__xor2_1 _09462_ (.A(_03063_),
    .B(_03064_),
    .X(_03066_));
 sky130_fd_sc_hd__inv_2 _09463_ (.A(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__and2_1 _09464_ (.A(_02901_),
    .B(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__xor2_1 _09465_ (.A(_02901_),
    .B(_03066_),
    .X(_03070_));
 sky130_fd_sc_hd__a21o_1 _09466_ (.A1(_02943_),
    .A2(_02952_),
    .B1(_02951_),
    .X(_03071_));
 sky130_fd_sc_hd__nand2_1 _09467_ (.A(_02914_),
    .B(_02918_),
    .Y(_03072_));
 sky130_fd_sc_hd__a31o_1 _09468_ (.A1(net7),
    .A2(net48),
    .A3(_02940_),
    .B1(_02939_),
    .X(_03073_));
 sky130_fd_sc_hd__nand4_2 _09469_ (.A(net6),
    .B(net7),
    .C(net49),
    .D(net50),
    .Y(_03074_));
 sky130_fd_sc_hd__a22o_1 _09470_ (.A1(net7),
    .A2(net49),
    .B1(net50),
    .B2(net6),
    .X(_03075_));
 sky130_fd_sc_hd__a22o_1 _09471_ (.A1(net5),
    .A2(net51),
    .B1(_03074_),
    .B2(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__nand4_2 _09472_ (.A(net5),
    .B(net51),
    .C(_03074_),
    .D(_03075_),
    .Y(_03077_));
 sky130_fd_sc_hd__nand3_2 _09473_ (.A(_03073_),
    .B(_03076_),
    .C(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__a21o_1 _09474_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_03073_),
    .X(_03079_));
 sky130_fd_sc_hd__nand3_2 _09475_ (.A(_03072_),
    .B(_03078_),
    .C(_03079_),
    .Y(_03081_));
 sky130_fd_sc_hd__a21o_1 _09476_ (.A1(_03078_),
    .A2(_03079_),
    .B1(_03072_),
    .X(_03082_));
 sky130_fd_sc_hd__and3_2 _09477_ (.A(_03071_),
    .B(_03081_),
    .C(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__a21oi_1 _09478_ (.A1(_03081_),
    .A2(_03082_),
    .B1(_03071_),
    .Y(_03084_));
 sky130_fd_sc_hd__a211oi_2 _09479_ (.A1(_02919_),
    .A2(_02921_),
    .B1(_03083_),
    .C1(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__a211o_1 _09480_ (.A1(_02919_),
    .A2(_02921_),
    .B1(_03083_),
    .C1(_03084_),
    .X(_03086_));
 sky130_fd_sc_hd__o211ai_1 _09481_ (.A1(_03083_),
    .A2(_03084_),
    .B1(_02919_),
    .C1(_02921_),
    .Y(_03087_));
 sky130_fd_sc_hd__o211a_1 _09482_ (.A1(_02923_),
    .A2(_02925_),
    .B1(_03086_),
    .C1(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__a211oi_1 _09483_ (.A1(_03086_),
    .A2(_03087_),
    .B1(_02923_),
    .C1(_02925_),
    .Y(_03089_));
 sky130_fd_sc_hd__or3_1 _09484_ (.A(_03070_),
    .B(_03088_),
    .C(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__o21ai_1 _09485_ (.A1(_03088_),
    .A2(_03089_),
    .B1(_03070_),
    .Y(_03092_));
 sky130_fd_sc_hd__o211a_2 _09486_ (.A1(_02974_),
    .A2(_02976_),
    .B1(_03090_),
    .C1(_03092_),
    .X(_03093_));
 sky130_fd_sc_hd__a211oi_2 _09487_ (.A1(_03090_),
    .A2(_03092_),
    .B1(_02974_),
    .C1(_02976_),
    .Y(_03094_));
 sky130_fd_sc_hd__a211oi_4 _09488_ (.A1(_02930_),
    .A2(_02932_),
    .B1(_03093_),
    .C1(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__o211a_1 _09489_ (.A1(_03093_),
    .A2(_03094_),
    .B1(_02930_),
    .C1(_02932_),
    .X(_03096_));
 sky130_fd_sc_hd__and4_1 _09490_ (.A(net9),
    .B(net10),
    .C(net46),
    .D(net47),
    .X(_03097_));
 sky130_fd_sc_hd__a22o_1 _09491_ (.A1(net10),
    .A2(net46),
    .B1(net47),
    .B2(net9),
    .X(_03098_));
 sky130_fd_sc_hd__and2b_1 _09492_ (.A_N(_03097_),
    .B(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__nand2_1 _09493_ (.A(net8),
    .B(net48),
    .Y(_03100_));
 sky130_fd_sc_hd__xnor2_2 _09494_ (.A(_03099_),
    .B(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__nand4_1 _09495_ (.A(net42),
    .B(net43),
    .C(net13),
    .D(net14),
    .Y(_03103_));
 sky130_fd_sc_hd__a22o_1 _09496_ (.A1(net43),
    .A2(net13),
    .B1(net14),
    .B2(net42),
    .X(_03104_));
 sky130_fd_sc_hd__and2_1 _09497_ (.A(net11),
    .B(net45),
    .X(_03105_));
 sky130_fd_sc_hd__a21o_1 _09498_ (.A1(_03103_),
    .A2(_03104_),
    .B1(_03105_),
    .X(_03106_));
 sky130_fd_sc_hd__nand3_1 _09499_ (.A(_03103_),
    .B(_03104_),
    .C(_03105_),
    .Y(_03107_));
 sky130_fd_sc_hd__a21bo_1 _09500_ (.A1(_02945_),
    .A2(_02946_),
    .B1_N(_02944_),
    .X(_03108_));
 sky130_fd_sc_hd__and3_1 _09501_ (.A(_03106_),
    .B(_03107_),
    .C(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__a21o_1 _09502_ (.A1(_03106_),
    .A2(_03107_),
    .B1(_03108_),
    .X(_03110_));
 sky130_fd_sc_hd__and2b_1 _09503_ (.A_N(_03109_),
    .B(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__xnor2_2 _09504_ (.A(_03101_),
    .B(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__nand2_1 _09505_ (.A(_02957_),
    .B(_02961_),
    .Y(_03114_));
 sky130_fd_sc_hd__a31o_1 _09506_ (.A1(net38),
    .A2(net17),
    .A3(_02981_),
    .B1(_02980_),
    .X(_03115_));
 sky130_fd_sc_hd__nand4_1 _09507_ (.A(net39),
    .B(net40),
    .C(net16),
    .D(net17),
    .Y(_03116_));
 sky130_fd_sc_hd__a22o_1 _09508_ (.A1(net40),
    .A2(net16),
    .B1(net17),
    .B2(net39),
    .X(_03117_));
 sky130_fd_sc_hd__a22o_1 _09509_ (.A1(net41),
    .A2(net15),
    .B1(_03116_),
    .B2(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__nand4_1 _09510_ (.A(net41),
    .B(net15),
    .C(_03116_),
    .D(_03117_),
    .Y(_03119_));
 sky130_fd_sc_hd__nand3_1 _09511_ (.A(_03115_),
    .B(_03118_),
    .C(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__a21o_1 _09512_ (.A1(_03118_),
    .A2(_03119_),
    .B1(_03115_),
    .X(_03121_));
 sky130_fd_sc_hd__nand3_1 _09513_ (.A(_03114_),
    .B(_03120_),
    .C(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__a21o_1 _09514_ (.A1(_03120_),
    .A2(_03121_),
    .B1(_03114_),
    .X(_03123_));
 sky130_fd_sc_hd__a21bo_1 _09515_ (.A1(_02955_),
    .A2(_02963_),
    .B1_N(_02962_),
    .X(_03125_));
 sky130_fd_sc_hd__and3_1 _09516_ (.A(_03122_),
    .B(_03123_),
    .C(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__inv_2 _09517_ (.A(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__a21oi_1 _09518_ (.A1(_03122_),
    .A2(_03123_),
    .B1(_03125_),
    .Y(_03128_));
 sky130_fd_sc_hd__nor3_1 _09519_ (.A(_03112_),
    .B(_03126_),
    .C(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__or3_2 _09520_ (.A(_03112_),
    .B(_03126_),
    .C(_03128_),
    .X(_03130_));
 sky130_fd_sc_hd__o21a_1 _09521_ (.A1(_03126_),
    .A2(_03128_),
    .B1(_03112_),
    .X(_03131_));
 sky130_fd_sc_hd__a211oi_4 _09522_ (.A1(_02997_),
    .A2(_02999_),
    .B1(_03129_),
    .C1(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__o211a_1 _09523_ (.A1(_03129_),
    .A2(_03131_),
    .B1(_02997_),
    .C1(_02999_),
    .X(_03133_));
 sky130_fd_sc_hd__a211oi_2 _09524_ (.A1(_02968_),
    .A2(_02972_),
    .B1(_03132_),
    .C1(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__o211a_1 _09525_ (.A1(_03132_),
    .A2(_03133_),
    .B1(_02968_),
    .C1(_02972_),
    .X(_03136_));
 sky130_fd_sc_hd__nand2_1 _09526_ (.A(_02992_),
    .B(_02995_),
    .Y(_03137_));
 sky130_fd_sc_hd__a21bo_1 _09527_ (.A1(_03001_),
    .A2(_03008_),
    .B1_N(_03007_),
    .X(_03138_));
 sky130_fd_sc_hd__and4_1 _09528_ (.A(net36),
    .B(net37),
    .C(net19),
    .D(net20),
    .X(_03139_));
 sky130_fd_sc_hd__a22o_1 _09529_ (.A1(net37),
    .A2(net19),
    .B1(net20),
    .B2(net36),
    .X(_03140_));
 sky130_fd_sc_hd__and2b_1 _09530_ (.A_N(_03139_),
    .B(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__nand2_1 _09531_ (.A(net38),
    .B(net18),
    .Y(_03142_));
 sky130_fd_sc_hd__xnor2_1 _09532_ (.A(_03141_),
    .B(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__nand4_1 _09533_ (.A(net64),
    .B(net34),
    .C(net22),
    .D(net24),
    .Y(_03144_));
 sky130_fd_sc_hd__a22o_1 _09534_ (.A1(net34),
    .A2(net22),
    .B1(net24),
    .B2(net64),
    .X(_03145_));
 sky130_fd_sc_hd__and2_1 _09535_ (.A(net35),
    .B(net21),
    .X(_03147_));
 sky130_fd_sc_hd__a21o_1 _09536_ (.A1(_03144_),
    .A2(_03145_),
    .B1(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__nand3_1 _09537_ (.A(_03144_),
    .B(_03145_),
    .C(_03147_),
    .Y(_03149_));
 sky130_fd_sc_hd__a21bo_1 _09538_ (.A1(_02987_),
    .A2(_02988_),
    .B1_N(_02986_),
    .X(_03150_));
 sky130_fd_sc_hd__nand3_1 _09539_ (.A(_03148_),
    .B(_03149_),
    .C(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__a21o_1 _09540_ (.A1(_03148_),
    .A2(_03149_),
    .B1(_03150_),
    .X(_03152_));
 sky130_fd_sc_hd__nand3_2 _09541_ (.A(_03143_),
    .B(_03151_),
    .C(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__a21o_1 _09542_ (.A1(_03151_),
    .A2(_03152_),
    .B1(_03143_),
    .X(_03154_));
 sky130_fd_sc_hd__nand3_4 _09543_ (.A(_03138_),
    .B(_03153_),
    .C(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__a21o_1 _09544_ (.A1(_03153_),
    .A2(_03154_),
    .B1(_03138_),
    .X(_03156_));
 sky130_fd_sc_hd__nand3_4 _09545_ (.A(_03137_),
    .B(_03155_),
    .C(_03156_),
    .Y(_03158_));
 sky130_fd_sc_hd__a21o_1 _09546_ (.A1(_03155_),
    .A2(_03156_),
    .B1(_03137_),
    .X(_03159_));
 sky130_fd_sc_hd__nand2_1 _09547_ (.A(_03002_),
    .B(_03006_),
    .Y(_03160_));
 sky130_fd_sc_hd__a22o_1 _09548_ (.A1(net63),
    .A2(net25),
    .B1(_03002_),
    .B2(_03003_),
    .X(_03161_));
 sky130_fd_sc_hd__nand4_2 _09549_ (.A(net63),
    .B(net25),
    .C(_03002_),
    .D(_03003_),
    .Y(_03162_));
 sky130_fd_sc_hd__nand3_2 _09550_ (.A(_02844_),
    .B(_03161_),
    .C(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__a21o_2 _09551_ (.A1(_03161_),
    .A2(_03162_),
    .B1(_02844_),
    .X(_03164_));
 sky130_fd_sc_hd__nand3_1 _09552_ (.A(_03160_),
    .B(_03163_),
    .C(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__a21o_1 _09553_ (.A1(_03163_),
    .A2(_03164_),
    .B1(_03160_),
    .X(_03166_));
 sky130_fd_sc_hd__nand3_1 _09554_ (.A(_02856_),
    .B(_03165_),
    .C(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__a21o_1 _09555_ (.A1(_03165_),
    .A2(_03166_),
    .B1(_02856_),
    .X(_03169_));
 sky130_fd_sc_hd__a31o_1 _09556_ (.A1(_02856_),
    .A2(_03009_),
    .A3(_03010_),
    .B1(_02854_),
    .X(_03170_));
 sky130_fd_sc_hd__nand3_4 _09557_ (.A(_03167_),
    .B(_03169_),
    .C(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__a21o_1 _09558_ (.A1(_03167_),
    .A2(_03169_),
    .B1(_03170_),
    .X(_03172_));
 sky130_fd_sc_hd__nand4_4 _09559_ (.A(_03158_),
    .B(_03159_),
    .C(_03171_),
    .D(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__a22o_1 _09560_ (.A1(_03158_),
    .A2(_03159_),
    .B1(_03171_),
    .B2(_03172_),
    .X(_03174_));
 sky130_fd_sc_hd__o211ai_4 _09561_ (.A1(_03016_),
    .A2(_03018_),
    .B1(_03173_),
    .C1(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__a211o_1 _09562_ (.A1(_03173_),
    .A2(_03174_),
    .B1(_03016_),
    .C1(_03018_),
    .X(_03176_));
 sky130_fd_sc_hd__or4bb_2 _09563_ (.A(_03134_),
    .B(_03136_),
    .C_N(_03175_),
    .D_N(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__a2bb2o_1 _09564_ (.A1_N(_03134_),
    .A2_N(_03136_),
    .B1(_03175_),
    .B2(_03176_),
    .X(_03178_));
 sky130_fd_sc_hd__o211a_2 _09565_ (.A1(_03021_),
    .A2(_03023_),
    .B1(_03177_),
    .C1(_03178_),
    .X(_03180_));
 sky130_fd_sc_hd__a211oi_2 _09566_ (.A1(_03177_),
    .A2(_03178_),
    .B1(_03021_),
    .C1(_03023_),
    .Y(_03181_));
 sky130_fd_sc_hd__nor4_2 _09567_ (.A(_03095_),
    .B(_03096_),
    .C(_03180_),
    .D(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__or4_1 _09568_ (.A(_03095_),
    .B(_03096_),
    .C(_03180_),
    .D(_03181_),
    .X(_03183_));
 sky130_fd_sc_hd__o22ai_1 _09569_ (.A1(_03095_),
    .A2(_03096_),
    .B1(_03180_),
    .B2(_03181_),
    .Y(_03184_));
 sky130_fd_sc_hd__o211a_1 _09570_ (.A1(_03025_),
    .A2(_03028_),
    .B1(_03183_),
    .C1(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__a211oi_1 _09571_ (.A1(_03183_),
    .A2(_03184_),
    .B1(_03025_),
    .C1(_03028_),
    .Y(_03186_));
 sky130_fd_sc_hd__nor2_1 _09572_ (.A(_03185_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__and2b_1 _09573_ (.A_N(_03050_),
    .B(_03187_),
    .X(_03188_));
 sky130_fd_sc_hd__xor2_2 _09574_ (.A(_03050_),
    .B(_03187_),
    .X(_03189_));
 sky130_fd_sc_hd__a21oi_2 _09575_ (.A1(_02891_),
    .A2(_03033_),
    .B1(_03032_),
    .Y(_03191_));
 sky130_fd_sc_hd__nor2_1 _09576_ (.A(_03189_),
    .B(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__xor2_2 _09577_ (.A(_03189_),
    .B(_03191_),
    .X(_03193_));
 sky130_fd_sc_hd__xnor2_2 _09578_ (.A(_03049_),
    .B(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__and2_1 _09579_ (.A(_03048_),
    .B(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__xnor2_1 _09580_ (.A(_03048_),
    .B(_03194_),
    .Y(_03196_));
 sky130_fd_sc_hd__a21bo_1 _09581_ (.A1(_03042_),
    .A2(_03046_),
    .B1_N(_03041_),
    .X(_03197_));
 sky130_fd_sc_hd__xnor2_1 _09582_ (.A(_03196_),
    .B(_03197_),
    .Y(net97));
 sky130_fd_sc_hd__nand2b_1 _09583_ (.A_N(_03088_),
    .B(_03090_),
    .Y(_03198_));
 sky130_fd_sc_hd__and4_1 _09584_ (.A(net4),
    .B(net5),
    .C(net52),
    .D(net53),
    .X(_03199_));
 sky130_fd_sc_hd__a22o_1 _09585_ (.A1(net5),
    .A2(net52),
    .B1(net53),
    .B2(net4),
    .X(_03201_));
 sky130_fd_sc_hd__and2b_1 _09586_ (.A_N(_03199_),
    .B(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__nand2_1 _09587_ (.A(net3),
    .B(net54),
    .Y(_03203_));
 sky130_fd_sc_hd__xnor2_1 _09588_ (.A(_03202_),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__a31o_1 _09589_ (.A1(net2),
    .A2(net54),
    .A3(_03052_),
    .B1(_03051_),
    .X(_03205_));
 sky130_fd_sc_hd__nand2_1 _09590_ (.A(_03204_),
    .B(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__xor2_1 _09591_ (.A(_03204_),
    .B(_03205_),
    .X(_03207_));
 sky130_fd_sc_hd__and4b_1 _09592_ (.A_N(net32),
    .B(net56),
    .C(net57),
    .D(net2),
    .X(_03208_));
 sky130_fd_sc_hd__o2bb2a_1 _09593_ (.A1_N(net2),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net32),
    .X(_03209_));
 sky130_fd_sc_hd__nor2_1 _09594_ (.A(_03208_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__xnor2_1 _09595_ (.A(_03207_),
    .B(_03210_),
    .Y(_03212_));
 sky130_fd_sc_hd__a21bo_1 _09596_ (.A1(_03059_),
    .A2(_03062_),
    .B1_N(_03057_),
    .X(_03213_));
 sky130_fd_sc_hd__nand2b_1 _09597_ (.A_N(_03212_),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__xor2_1 _09598_ (.A(_03212_),
    .B(_03213_),
    .X(_03215_));
 sky130_fd_sc_hd__inv_2 _09599_ (.A(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__nand2_1 _09600_ (.A(_03060_),
    .B(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__xor2_1 _09601_ (.A(_03060_),
    .B(_03215_),
    .X(_03218_));
 sky130_fd_sc_hd__a21o_1 _09602_ (.A1(_03101_),
    .A2(_03110_),
    .B1(_03109_),
    .X(_03219_));
 sky130_fd_sc_hd__nand2_1 _09603_ (.A(_03074_),
    .B(_03077_),
    .Y(_03220_));
 sky130_fd_sc_hd__a31o_1 _09604_ (.A1(net8),
    .A2(net48),
    .A3(_03098_),
    .B1(_03097_),
    .X(_03221_));
 sky130_fd_sc_hd__nand4_2 _09605_ (.A(net7),
    .B(net8),
    .C(net49),
    .D(net50),
    .Y(_03223_));
 sky130_fd_sc_hd__a22o_1 _09606_ (.A1(net8),
    .A2(net49),
    .B1(net50),
    .B2(net7),
    .X(_03224_));
 sky130_fd_sc_hd__a22o_1 _09607_ (.A1(net6),
    .A2(net51),
    .B1(_03223_),
    .B2(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__nand4_2 _09608_ (.A(net6),
    .B(net51),
    .C(_03223_),
    .D(_03224_),
    .Y(_03226_));
 sky130_fd_sc_hd__nand3_2 _09609_ (.A(_03221_),
    .B(_03225_),
    .C(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__a21o_1 _09610_ (.A1(_03225_),
    .A2(_03226_),
    .B1(_03221_),
    .X(_03228_));
 sky130_fd_sc_hd__nand3_2 _09611_ (.A(_03220_),
    .B(_03227_),
    .C(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__a21o_1 _09612_ (.A1(_03227_),
    .A2(_03228_),
    .B1(_03220_),
    .X(_03230_));
 sky130_fd_sc_hd__and3_1 _09613_ (.A(_03219_),
    .B(_03229_),
    .C(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__nand3_1 _09614_ (.A(_03219_),
    .B(_03229_),
    .C(_03230_),
    .Y(_03232_));
 sky130_fd_sc_hd__a21oi_1 _09615_ (.A1(_03229_),
    .A2(_03230_),
    .B1(_03219_),
    .Y(_03234_));
 sky130_fd_sc_hd__a211o_1 _09616_ (.A1(_03078_),
    .A2(_03081_),
    .B1(_03231_),
    .C1(_03234_),
    .X(_03235_));
 sky130_fd_sc_hd__o211ai_2 _09617_ (.A1(_03231_),
    .A2(_03234_),
    .B1(_03078_),
    .C1(_03081_),
    .Y(_03236_));
 sky130_fd_sc_hd__o211a_2 _09618_ (.A1(_03083_),
    .A2(_03085_),
    .B1(_03235_),
    .C1(_03236_),
    .X(_03237_));
 sky130_fd_sc_hd__a211oi_2 _09619_ (.A1(_03235_),
    .A2(_03236_),
    .B1(_03083_),
    .C1(_03085_),
    .Y(_03238_));
 sky130_fd_sc_hd__nor3_1 _09620_ (.A(_03218_),
    .B(_03237_),
    .C(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__or3_2 _09621_ (.A(_03218_),
    .B(_03237_),
    .C(_03238_),
    .X(_03240_));
 sky130_fd_sc_hd__o21ai_2 _09622_ (.A1(_03237_),
    .A2(_03238_),
    .B1(_03218_),
    .Y(_03241_));
 sky130_fd_sc_hd__o211ai_4 _09623_ (.A1(_03132_),
    .A2(_03134_),
    .B1(_03240_),
    .C1(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__a211o_1 _09624_ (.A1(_03240_),
    .A2(_03241_),
    .B1(_03132_),
    .C1(_03134_),
    .X(_03243_));
 sky130_fd_sc_hd__nand3_4 _09625_ (.A(_03198_),
    .B(_03242_),
    .C(_03243_),
    .Y(_03245_));
 sky130_fd_sc_hd__a21o_1 _09626_ (.A1(_03242_),
    .A2(_03243_),
    .B1(_03198_),
    .X(_03246_));
 sky130_fd_sc_hd__and4_1 _09627_ (.A(net10),
    .B(net11),
    .C(net46),
    .D(net47),
    .X(_03247_));
 sky130_fd_sc_hd__a22o_1 _09628_ (.A1(net11),
    .A2(net46),
    .B1(net47),
    .B2(net10),
    .X(_03248_));
 sky130_fd_sc_hd__and2b_1 _09629_ (.A_N(_03247_),
    .B(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__nand2_1 _09630_ (.A(net9),
    .B(net48),
    .Y(_03250_));
 sky130_fd_sc_hd__xnor2_2 _09631_ (.A(_03249_),
    .B(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__nand4_1 _09632_ (.A(net42),
    .B(net43),
    .C(net14),
    .D(net15),
    .Y(_03252_));
 sky130_fd_sc_hd__a22o_1 _09633_ (.A1(net43),
    .A2(net14),
    .B1(net15),
    .B2(net42),
    .X(_03253_));
 sky130_fd_sc_hd__and2_1 _09634_ (.A(net13),
    .B(net45),
    .X(_03254_));
 sky130_fd_sc_hd__a21o_1 _09635_ (.A1(_03252_),
    .A2(_03253_),
    .B1(_03254_),
    .X(_03256_));
 sky130_fd_sc_hd__nand3_1 _09636_ (.A(_03252_),
    .B(_03253_),
    .C(_03254_),
    .Y(_03257_));
 sky130_fd_sc_hd__a21bo_1 _09637_ (.A1(_03104_),
    .A2(_03105_),
    .B1_N(_03103_),
    .X(_03258_));
 sky130_fd_sc_hd__and3_1 _09638_ (.A(_03256_),
    .B(_03257_),
    .C(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__a21o_1 _09639_ (.A1(_03256_),
    .A2(_03257_),
    .B1(_03258_),
    .X(_03260_));
 sky130_fd_sc_hd__and2b_1 _09640_ (.A_N(_03259_),
    .B(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__xnor2_2 _09641_ (.A(_03251_),
    .B(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _09642_ (.A(_03116_),
    .B(_03119_),
    .Y(_03263_));
 sky130_fd_sc_hd__a31o_1 _09643_ (.A1(net38),
    .A2(net18),
    .A3(_03140_),
    .B1(_03139_),
    .X(_03264_));
 sky130_fd_sc_hd__nand4_1 _09644_ (.A(net39),
    .B(net40),
    .C(net17),
    .D(net18),
    .Y(_03265_));
 sky130_fd_sc_hd__a22o_1 _09645_ (.A1(net40),
    .A2(net17),
    .B1(net18),
    .B2(net39),
    .X(_03267_));
 sky130_fd_sc_hd__a22o_1 _09646_ (.A1(net41),
    .A2(net16),
    .B1(_03265_),
    .B2(_03267_),
    .X(_03268_));
 sky130_fd_sc_hd__nand4_1 _09647_ (.A(net41),
    .B(net16),
    .C(_03265_),
    .D(_03267_),
    .Y(_03269_));
 sky130_fd_sc_hd__nand3_1 _09648_ (.A(_03264_),
    .B(_03268_),
    .C(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__a21o_1 _09649_ (.A1(_03268_),
    .A2(_03269_),
    .B1(_03264_),
    .X(_03271_));
 sky130_fd_sc_hd__nand3_1 _09650_ (.A(_03263_),
    .B(_03270_),
    .C(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__a21o_1 _09651_ (.A1(_03270_),
    .A2(_03271_),
    .B1(_03263_),
    .X(_03273_));
 sky130_fd_sc_hd__a21bo_1 _09652_ (.A1(_03114_),
    .A2(_03121_),
    .B1_N(_03120_),
    .X(_03274_));
 sky130_fd_sc_hd__and3_1 _09653_ (.A(_03272_),
    .B(_03273_),
    .C(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__inv_2 _09654_ (.A(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__a21oi_1 _09655_ (.A1(_03272_),
    .A2(_03273_),
    .B1(_03274_),
    .Y(_03278_));
 sky130_fd_sc_hd__nor3_2 _09656_ (.A(_03262_),
    .B(_03275_),
    .C(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__inv_2 _09657_ (.A(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__o21a_1 _09658_ (.A1(_03275_),
    .A2(_03278_),
    .B1(_03262_),
    .X(_03281_));
 sky130_fd_sc_hd__a211oi_4 _09659_ (.A1(_03155_),
    .A2(_03158_),
    .B1(_03279_),
    .C1(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__o211a_1 _09660_ (.A1(_03279_),
    .A2(_03281_),
    .B1(_03155_),
    .C1(_03158_),
    .X(_03283_));
 sky130_fd_sc_hd__a211oi_4 _09661_ (.A1(_03127_),
    .A2(_03130_),
    .B1(_03282_),
    .C1(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__o211a_1 _09662_ (.A1(_03282_),
    .A2(_03283_),
    .B1(_03127_),
    .C1(_03130_),
    .X(_03285_));
 sky130_fd_sc_hd__nand2_1 _09663_ (.A(_03151_),
    .B(_03153_),
    .Y(_03286_));
 sky130_fd_sc_hd__a21bo_1 _09664_ (.A1(_03160_),
    .A2(_03164_),
    .B1_N(_03163_),
    .X(_03287_));
 sky130_fd_sc_hd__and4_1 _09665_ (.A(net36),
    .B(net37),
    .C(net20),
    .D(net21),
    .X(_03289_));
 sky130_fd_sc_hd__a22o_1 _09666_ (.A1(net37),
    .A2(net20),
    .B1(net21),
    .B2(net36),
    .X(_03290_));
 sky130_fd_sc_hd__and2b_1 _09667_ (.A_N(_03289_),
    .B(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__nand2_1 _09668_ (.A(net38),
    .B(net19),
    .Y(_03292_));
 sky130_fd_sc_hd__xnor2_1 _09669_ (.A(_03291_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__and3_1 _09670_ (.A(net64),
    .B(net34),
    .C(net25),
    .X(_03294_));
 sky130_fd_sc_hd__nand4_1 _09671_ (.A(net64),
    .B(net34),
    .C(net24),
    .D(net25),
    .Y(_03295_));
 sky130_fd_sc_hd__a22o_1 _09672_ (.A1(net34),
    .A2(net24),
    .B1(net25),
    .B2(net64),
    .X(_03296_));
 sky130_fd_sc_hd__and2_1 _09673_ (.A(net35),
    .B(net22),
    .X(_03297_));
 sky130_fd_sc_hd__a21o_1 _09674_ (.A1(_03295_),
    .A2(_03296_),
    .B1(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__nand3_1 _09675_ (.A(_03295_),
    .B(_03296_),
    .C(_03297_),
    .Y(_03300_));
 sky130_fd_sc_hd__a21bo_1 _09676_ (.A1(_03145_),
    .A2(_03147_),
    .B1_N(_03144_),
    .X(_03301_));
 sky130_fd_sc_hd__nand3_1 _09677_ (.A(_03298_),
    .B(_03300_),
    .C(_03301_),
    .Y(_03302_));
 sky130_fd_sc_hd__a21o_1 _09678_ (.A1(_03298_),
    .A2(_03300_),
    .B1(_03301_),
    .X(_03303_));
 sky130_fd_sc_hd__nand3_2 _09679_ (.A(_03293_),
    .B(_03302_),
    .C(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__a21o_1 _09680_ (.A1(_03302_),
    .A2(_03303_),
    .B1(_03293_),
    .X(_03305_));
 sky130_fd_sc_hd__nand3_4 _09681_ (.A(_03287_),
    .B(_03304_),
    .C(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__a21o_1 _09682_ (.A1(_03304_),
    .A2(_03305_),
    .B1(_03287_),
    .X(_03307_));
 sky130_fd_sc_hd__nand3_4 _09683_ (.A(_03286_),
    .B(_03306_),
    .C(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__a21o_1 _09684_ (.A1(_03306_),
    .A2(_03307_),
    .B1(_03286_),
    .X(_03309_));
 sky130_fd_sc_hd__a31oi_2 _09685_ (.A1(_02856_),
    .A2(_03165_),
    .A3(_03166_),
    .B1(_02854_),
    .Y(_03311_));
 sky130_fd_sc_hd__nand2_2 _09686_ (.A(_03002_),
    .B(_03162_),
    .Y(_03312_));
 sky130_fd_sc_hd__nand3_1 _09687_ (.A(_03163_),
    .B(_03164_),
    .C(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__a21o_1 _09688_ (.A1(_03163_),
    .A2(_03164_),
    .B1(_03312_),
    .X(_03314_));
 sky130_fd_sc_hd__nand2_1 _09689_ (.A(_03313_),
    .B(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__a21bo_1 _09690_ (.A1(_03313_),
    .A2(_03314_),
    .B1_N(_02856_),
    .X(_03316_));
 sky130_fd_sc_hd__nand3b_1 _09691_ (.A_N(_02856_),
    .B(_03313_),
    .C(_03314_),
    .Y(_03317_));
 sky130_fd_sc_hd__a21oi_1 _09692_ (.A1(_03316_),
    .A2(_03317_),
    .B1(_03311_),
    .Y(_03318_));
 sky130_fd_sc_hd__a21o_1 _09693_ (.A1(_03316_),
    .A2(_03317_),
    .B1(_03311_),
    .X(_03319_));
 sky130_fd_sc_hd__nand3_2 _09694_ (.A(_03311_),
    .B(_03316_),
    .C(_03317_),
    .Y(_03320_));
 sky130_fd_sc_hd__and4_1 _09695_ (.A(_03308_),
    .B(_03309_),
    .C(_03319_),
    .D(_03320_),
    .X(_03322_));
 sky130_fd_sc_hd__a22oi_4 _09696_ (.A1(_03308_),
    .A2(_03309_),
    .B1(_03319_),
    .B2(_03320_),
    .Y(_03323_));
 sky130_fd_sc_hd__a211oi_4 _09697_ (.A1(_03171_),
    .A2(_03173_),
    .B1(_03322_),
    .C1(_03323_),
    .Y(_03324_));
 sky130_fd_sc_hd__o211a_1 _09698_ (.A1(_03322_),
    .A2(_03323_),
    .B1(_03171_),
    .C1(_03173_),
    .X(_03325_));
 sky130_fd_sc_hd__nor4_2 _09699_ (.A(_03284_),
    .B(_03285_),
    .C(_03324_),
    .D(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__o22a_1 _09700_ (.A1(_03284_),
    .A2(_03285_),
    .B1(_03324_),
    .B2(_03325_),
    .X(_03327_));
 sky130_fd_sc_hd__a211o_2 _09701_ (.A1(_03175_),
    .A2(_03177_),
    .B1(_03326_),
    .C1(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__o211ai_2 _09702_ (.A1(_03326_),
    .A2(_03327_),
    .B1(_03175_),
    .C1(_03177_),
    .Y(_03329_));
 sky130_fd_sc_hd__nand4_4 _09703_ (.A(_03245_),
    .B(_03246_),
    .C(_03328_),
    .D(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__a22o_1 _09704_ (.A1(_03245_),
    .A2(_03246_),
    .B1(_03328_),
    .B2(_03329_),
    .X(_03331_));
 sky130_fd_sc_hd__o211ai_4 _09705_ (.A1(_03180_),
    .A2(_03182_),
    .B1(_03330_),
    .C1(_03331_),
    .Y(_03333_));
 sky130_fd_sc_hd__a211o_1 _09706_ (.A1(_03330_),
    .A2(_03331_),
    .B1(_03180_),
    .C1(_03182_),
    .X(_03334_));
 sky130_fd_sc_hd__o211ai_4 _09707_ (.A1(_03093_),
    .A2(_03095_),
    .B1(_03333_),
    .C1(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__a211o_1 _09708_ (.A1(_03333_),
    .A2(_03334_),
    .B1(_03093_),
    .C1(_03095_),
    .X(_03336_));
 sky130_fd_sc_hd__o211ai_4 _09709_ (.A1(_03185_),
    .A2(_03188_),
    .B1(_03335_),
    .C1(_03336_),
    .Y(_03337_));
 sky130_fd_sc_hd__a211o_1 _09710_ (.A1(_03335_),
    .A2(_03336_),
    .B1(_03185_),
    .C1(_03188_),
    .X(_03338_));
 sky130_fd_sc_hd__o211ai_4 _09711_ (.A1(_03065_),
    .A2(_03068_),
    .B1(_03337_),
    .C1(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__a211o_1 _09712_ (.A1(_03337_),
    .A2(_03338_),
    .B1(_03065_),
    .C1(_03068_),
    .X(_03340_));
 sky130_fd_sc_hd__nand2_1 _09713_ (.A(_03339_),
    .B(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__a21o_1 _09714_ (.A1(_03049_),
    .A2(_03193_),
    .B1(_03192_),
    .X(_03342_));
 sky130_fd_sc_hd__xor2_1 _09715_ (.A(_03341_),
    .B(_03342_),
    .X(_03344_));
 sky130_fd_sc_hd__nor2_1 _09716_ (.A(_03043_),
    .B(_03196_),
    .Y(_03345_));
 sky130_fd_sc_hd__o21a_1 _09717_ (.A1(_03048_),
    .A2(_03194_),
    .B1(_03041_),
    .X(_03346_));
 sky130_fd_sc_hd__a2bb2o_1 _09718_ (.A1_N(_03195_),
    .A2_N(_03346_),
    .B1(_03345_),
    .B2(_03044_),
    .X(_03347_));
 sky130_fd_sc_hd__a31oi_4 _09719_ (.A1(_02727_),
    .A2(_03045_),
    .A3(_03345_),
    .B1(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__and4_1 _09720_ (.A(_02390_),
    .B(_02725_),
    .C(_03045_),
    .D(_03345_),
    .X(_03349_));
 sky130_fd_sc_hd__o31ai_4 _09721_ (.A1(_02049_),
    .A2(_02051_),
    .A3(_02052_),
    .B1(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__and2_1 _09722_ (.A(_03348_),
    .B(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__a21oi_1 _09723_ (.A1(_03348_),
    .A2(_03350_),
    .B1(_03344_),
    .Y(_03352_));
 sky130_fd_sc_hd__and3_1 _09724_ (.A(_03344_),
    .B(_03348_),
    .C(_03350_),
    .X(_03353_));
 sky130_fd_sc_hd__nor2_1 _09725_ (.A(_03352_),
    .B(_03353_),
    .Y(net99));
 sky130_fd_sc_hd__and4_1 _09726_ (.A(net5),
    .B(net6),
    .C(net52),
    .D(net53),
    .X(_03355_));
 sky130_fd_sc_hd__a22o_1 _09727_ (.A1(net6),
    .A2(net52),
    .B1(net53),
    .B2(net5),
    .X(_03356_));
 sky130_fd_sc_hd__and2b_1 _09728_ (.A_N(_03355_),
    .B(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__nand2_1 _09729_ (.A(net4),
    .B(net54),
    .Y(_03358_));
 sky130_fd_sc_hd__xnor2_1 _09730_ (.A(_03357_),
    .B(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__a31o_1 _09731_ (.A1(net3),
    .A2(net54),
    .A3(_03201_),
    .B1(_03199_),
    .X(_03360_));
 sky130_fd_sc_hd__nand2_1 _09732_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__xor2_1 _09733_ (.A(_03359_),
    .B(_03360_),
    .X(_03362_));
 sky130_fd_sc_hd__and4b_1 _09734_ (.A_N(net2),
    .B(net3),
    .C(net56),
    .D(net57),
    .X(_03363_));
 sky130_fd_sc_hd__o2bb2a_1 _09735_ (.A1_N(net3),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net2),
    .X(_03364_));
 sky130_fd_sc_hd__nor2_1 _09736_ (.A(_03363_),
    .B(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__xnor2_1 _09737_ (.A(_03362_),
    .B(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__a21bo_1 _09738_ (.A1(_03207_),
    .A2(_03210_),
    .B1_N(_03206_),
    .X(_03367_));
 sky130_fd_sc_hd__and2b_1 _09739_ (.A_N(_03366_),
    .B(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__xor2_1 _09740_ (.A(_03366_),
    .B(_03367_),
    .X(_03369_));
 sky130_fd_sc_hd__inv_2 _09741_ (.A(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__and2_1 _09742_ (.A(_03208_),
    .B(_03370_),
    .X(_03371_));
 sky130_fd_sc_hd__xor2_1 _09743_ (.A(_03208_),
    .B(_03369_),
    .X(_03372_));
 sky130_fd_sc_hd__a21o_1 _09744_ (.A1(_03251_),
    .A2(_03260_),
    .B1(_03259_),
    .X(_03373_));
 sky130_fd_sc_hd__nand2_1 _09745_ (.A(_03223_),
    .B(_03226_),
    .Y(_03375_));
 sky130_fd_sc_hd__a31o_1 _09746_ (.A1(net9),
    .A2(net48),
    .A3(_03248_),
    .B1(_03247_),
    .X(_03376_));
 sky130_fd_sc_hd__nand4_2 _09747_ (.A(net8),
    .B(net9),
    .C(net49),
    .D(net50),
    .Y(_03377_));
 sky130_fd_sc_hd__a22o_1 _09748_ (.A1(net9),
    .A2(net49),
    .B1(net50),
    .B2(net8),
    .X(_03378_));
 sky130_fd_sc_hd__a22o_1 _09749_ (.A1(net7),
    .A2(net51),
    .B1(_03377_),
    .B2(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__nand4_2 _09750_ (.A(net7),
    .B(net51),
    .C(_03377_),
    .D(_03378_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand3_2 _09751_ (.A(_03376_),
    .B(_03379_),
    .C(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__a21o_1 _09752_ (.A1(_03379_),
    .A2(_03380_),
    .B1(_03376_),
    .X(_03382_));
 sky130_fd_sc_hd__nand3_1 _09753_ (.A(_03375_),
    .B(_03381_),
    .C(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__a21o_1 _09754_ (.A1(_03381_),
    .A2(_03382_),
    .B1(_03375_),
    .X(_03384_));
 sky130_fd_sc_hd__and3_1 _09755_ (.A(_03373_),
    .B(_03383_),
    .C(_03384_),
    .X(_03386_));
 sky130_fd_sc_hd__a21oi_1 _09756_ (.A1(_03383_),
    .A2(_03384_),
    .B1(_03373_),
    .Y(_03387_));
 sky130_fd_sc_hd__a211oi_2 _09757_ (.A1(_03227_),
    .A2(_03229_),
    .B1(_03386_),
    .C1(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__o211a_1 _09758_ (.A1(_03386_),
    .A2(_03387_),
    .B1(_03227_),
    .C1(_03229_),
    .X(_03389_));
 sky130_fd_sc_hd__a211oi_2 _09759_ (.A1(_03232_),
    .A2(_03235_),
    .B1(_03388_),
    .C1(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__o211a_1 _09760_ (.A1(_03388_),
    .A2(_03389_),
    .B1(_03232_),
    .C1(_03235_),
    .X(_03391_));
 sky130_fd_sc_hd__or3_2 _09761_ (.A(_03372_),
    .B(_03390_),
    .C(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__o21ai_2 _09762_ (.A1(_03390_),
    .A2(_03391_),
    .B1(_03372_),
    .Y(_03393_));
 sky130_fd_sc_hd__o211a_1 _09763_ (.A1(_03282_),
    .A2(_03284_),
    .B1(_03392_),
    .C1(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__o211ai_2 _09764_ (.A1(_03282_),
    .A2(_03284_),
    .B1(_03392_),
    .C1(_03393_),
    .Y(_03395_));
 sky130_fd_sc_hd__a211o_1 _09765_ (.A1(_03392_),
    .A2(_03393_),
    .B1(_03282_),
    .C1(_03284_),
    .X(_03397_));
 sky130_fd_sc_hd__o211a_2 _09766_ (.A1(_03237_),
    .A2(_03239_),
    .B1(_03395_),
    .C1(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__a211oi_2 _09767_ (.A1(_03395_),
    .A2(_03397_),
    .B1(_03237_),
    .C1(_03239_),
    .Y(_03399_));
 sky130_fd_sc_hd__and4_1 _09768_ (.A(net11),
    .B(net13),
    .C(net46),
    .D(net47),
    .X(_03400_));
 sky130_fd_sc_hd__a22o_1 _09769_ (.A1(net13),
    .A2(net46),
    .B1(net47),
    .B2(net11),
    .X(_03401_));
 sky130_fd_sc_hd__and2b_1 _09770_ (.A_N(_03400_),
    .B(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__nand2_1 _09771_ (.A(net10),
    .B(net48),
    .Y(_03403_));
 sky130_fd_sc_hd__xnor2_2 _09772_ (.A(_03402_),
    .B(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand4_1 _09773_ (.A(net42),
    .B(net43),
    .C(net15),
    .D(net16),
    .Y(_03405_));
 sky130_fd_sc_hd__a22o_1 _09774_ (.A1(net43),
    .A2(net15),
    .B1(net16),
    .B2(net42),
    .X(_03406_));
 sky130_fd_sc_hd__and2_1 _09775_ (.A(net45),
    .B(net14),
    .X(_03408_));
 sky130_fd_sc_hd__a21o_1 _09776_ (.A1(_03405_),
    .A2(_03406_),
    .B1(_03408_),
    .X(_03409_));
 sky130_fd_sc_hd__nand3_1 _09777_ (.A(_03405_),
    .B(_03406_),
    .C(_03408_),
    .Y(_03410_));
 sky130_fd_sc_hd__a21bo_1 _09778_ (.A1(_03253_),
    .A2(_03254_),
    .B1_N(_03252_),
    .X(_03411_));
 sky130_fd_sc_hd__and3_1 _09779_ (.A(_03409_),
    .B(_03410_),
    .C(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__a21o_1 _09780_ (.A1(_03409_),
    .A2(_03410_),
    .B1(_03411_),
    .X(_03413_));
 sky130_fd_sc_hd__and2b_1 _09781_ (.A_N(_03412_),
    .B(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__xnor2_2 _09782_ (.A(_03404_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand2_1 _09783_ (.A(_03265_),
    .B(_03269_),
    .Y(_03416_));
 sky130_fd_sc_hd__a31o_1 _09784_ (.A1(net38),
    .A2(net19),
    .A3(_03290_),
    .B1(_03289_),
    .X(_03417_));
 sky130_fd_sc_hd__nand4_1 _09785_ (.A(net39),
    .B(net40),
    .C(net18),
    .D(net19),
    .Y(_03419_));
 sky130_fd_sc_hd__a22o_1 _09786_ (.A1(net40),
    .A2(net18),
    .B1(net19),
    .B2(net39),
    .X(_03420_));
 sky130_fd_sc_hd__a22o_1 _09787_ (.A1(net41),
    .A2(net17),
    .B1(_03419_),
    .B2(_03420_),
    .X(_03421_));
 sky130_fd_sc_hd__nand4_1 _09788_ (.A(net41),
    .B(net17),
    .C(_03419_),
    .D(_03420_),
    .Y(_03422_));
 sky130_fd_sc_hd__nand3_1 _09789_ (.A(_03417_),
    .B(_03421_),
    .C(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21o_1 _09790_ (.A1(_03421_),
    .A2(_03422_),
    .B1(_03417_),
    .X(_03424_));
 sky130_fd_sc_hd__nand3_1 _09791_ (.A(_03416_),
    .B(_03423_),
    .C(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__a21o_1 _09792_ (.A1(_03423_),
    .A2(_03424_),
    .B1(_03416_),
    .X(_03426_));
 sky130_fd_sc_hd__a21bo_1 _09793_ (.A1(_03263_),
    .A2(_03271_),
    .B1_N(_03270_),
    .X(_03427_));
 sky130_fd_sc_hd__and3_1 _09794_ (.A(_03425_),
    .B(_03426_),
    .C(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__inv_2 _09795_ (.A(_03428_),
    .Y(_03430_));
 sky130_fd_sc_hd__a21oi_1 _09796_ (.A1(_03425_),
    .A2(_03426_),
    .B1(_03427_),
    .Y(_03431_));
 sky130_fd_sc_hd__nor3_1 _09797_ (.A(_03415_),
    .B(_03428_),
    .C(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__or3_1 _09798_ (.A(_03415_),
    .B(_03428_),
    .C(_03431_),
    .X(_03433_));
 sky130_fd_sc_hd__o21a_1 _09799_ (.A1(_03428_),
    .A2(_03431_),
    .B1(_03415_),
    .X(_03434_));
 sky130_fd_sc_hd__a211oi_4 _09800_ (.A1(_03306_),
    .A2(_03308_),
    .B1(_03432_),
    .C1(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__o211a_1 _09801_ (.A1(_03432_),
    .A2(_03434_),
    .B1(_03306_),
    .C1(_03308_),
    .X(_03436_));
 sky130_fd_sc_hd__a211oi_4 _09802_ (.A1(_03276_),
    .A2(_03280_),
    .B1(_03435_),
    .C1(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__o211a_1 _09803_ (.A1(_03435_),
    .A2(_03436_),
    .B1(_03276_),
    .C1(_03280_),
    .X(_03438_));
 sky130_fd_sc_hd__nand2_1 _09804_ (.A(_03302_),
    .B(_03304_),
    .Y(_03439_));
 sky130_fd_sc_hd__a21boi_4 _09805_ (.A1(_03164_),
    .A2(_03312_),
    .B1_N(_03163_),
    .Y(_03441_));
 sky130_fd_sc_hd__a21bo_1 _09806_ (.A1(_03164_),
    .A2(_03312_),
    .B1_N(_03163_),
    .X(_03442_));
 sky130_fd_sc_hd__and4_1 _09807_ (.A(net36),
    .B(net37),
    .C(net21),
    .D(net22),
    .X(_03443_));
 sky130_fd_sc_hd__a22o_1 _09808_ (.A1(net37),
    .A2(net21),
    .B1(net22),
    .B2(net36),
    .X(_03444_));
 sky130_fd_sc_hd__and2b_1 _09809_ (.A_N(_03443_),
    .B(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__nand2_1 _09810_ (.A(net38),
    .B(net20),
    .Y(_03446_));
 sky130_fd_sc_hd__xnor2_1 _09811_ (.A(_03445_),
    .B(_03446_),
    .Y(_03447_));
 sky130_fd_sc_hd__o21ai_2 _09812_ (.A1(net64),
    .A2(net34),
    .B1(net25),
    .Y(_03448_));
 sky130_fd_sc_hd__nand2_1 _09813_ (.A(net35),
    .B(net24),
    .Y(_03449_));
 sky130_fd_sc_hd__o21ai_1 _09814_ (.A1(_03294_),
    .A2(_03448_),
    .B1(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__or3_1 _09815_ (.A(_03294_),
    .B(_03448_),
    .C(_03449_),
    .X(_03452_));
 sky130_fd_sc_hd__a21bo_1 _09816_ (.A1(_03296_),
    .A2(_03297_),
    .B1_N(_03295_),
    .X(_03453_));
 sky130_fd_sc_hd__nand3_1 _09817_ (.A(_03450_),
    .B(_03452_),
    .C(_03453_),
    .Y(_03454_));
 sky130_fd_sc_hd__a21o_1 _09818_ (.A1(_03450_),
    .A2(_03452_),
    .B1(_03453_),
    .X(_03455_));
 sky130_fd_sc_hd__nand3_1 _09819_ (.A(_03447_),
    .B(_03454_),
    .C(_03455_),
    .Y(_03456_));
 sky130_fd_sc_hd__a21o_1 _09820_ (.A1(_03454_),
    .A2(_03455_),
    .B1(_03447_),
    .X(_03457_));
 sky130_fd_sc_hd__nand3_2 _09821_ (.A(_03442_),
    .B(_03456_),
    .C(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__a21o_1 _09822_ (.A1(_03456_),
    .A2(_03457_),
    .B1(_03442_),
    .X(_03459_));
 sky130_fd_sc_hd__nand3_2 _09823_ (.A(_03439_),
    .B(_03458_),
    .C(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__a21o_1 _09824_ (.A1(_03458_),
    .A2(_03459_),
    .B1(_03439_),
    .X(_03461_));
 sky130_fd_sc_hd__and3_4 _09825_ (.A(_02854_),
    .B(_03313_),
    .C(_03314_),
    .X(_03463_));
 sky130_fd_sc_hd__inv_2 _09826_ (.A(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__a21oi_4 _09827_ (.A1(_02855_),
    .A2(_03315_),
    .B1(_03463_),
    .Y(_03465_));
 sky130_fd_sc_hd__a21o_1 _09828_ (.A1(_02855_),
    .A2(_03315_),
    .B1(_03463_),
    .X(_03466_));
 sky130_fd_sc_hd__nand3_1 _09829_ (.A(_03460_),
    .B(_03461_),
    .C(_03465_),
    .Y(_03467_));
 sky130_fd_sc_hd__a21o_1 _09830_ (.A1(_03460_),
    .A2(_03461_),
    .B1(_03465_),
    .X(_03468_));
 sky130_fd_sc_hd__a31o_1 _09831_ (.A1(_03308_),
    .A2(_03309_),
    .A3(_03320_),
    .B1(_03318_),
    .X(_03469_));
 sky130_fd_sc_hd__and3_2 _09832_ (.A(_03467_),
    .B(_03468_),
    .C(_03469_),
    .X(_03470_));
 sky130_fd_sc_hd__a21oi_2 _09833_ (.A1(_03467_),
    .A2(_03468_),
    .B1(_03469_),
    .Y(_03471_));
 sky130_fd_sc_hd__nor4_2 _09834_ (.A(_03437_),
    .B(_03438_),
    .C(_03470_),
    .D(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__or4_1 _09835_ (.A(_03437_),
    .B(_03438_),
    .C(_03470_),
    .D(_03471_),
    .X(_03474_));
 sky130_fd_sc_hd__o22ai_2 _09836_ (.A1(_03437_),
    .A2(_03438_),
    .B1(_03470_),
    .B2(_03471_),
    .Y(_03475_));
 sky130_fd_sc_hd__o211a_2 _09837_ (.A1(_03324_),
    .A2(_03326_),
    .B1(_03474_),
    .C1(_03475_),
    .X(_03476_));
 sky130_fd_sc_hd__a211oi_2 _09838_ (.A1(_03474_),
    .A2(_03475_),
    .B1(_03324_),
    .C1(_03326_),
    .Y(_03477_));
 sky130_fd_sc_hd__nor4_4 _09839_ (.A(_03398_),
    .B(_03399_),
    .C(_03476_),
    .D(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__o22a_1 _09840_ (.A1(_03398_),
    .A2(_03399_),
    .B1(_03476_),
    .B2(_03477_),
    .X(_03479_));
 sky130_fd_sc_hd__a211oi_4 _09841_ (.A1(_03328_),
    .A2(_03330_),
    .B1(_03478_),
    .C1(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__o211a_1 _09842_ (.A1(_03478_),
    .A2(_03479_),
    .B1(_03328_),
    .C1(_03330_),
    .X(_03481_));
 sky130_fd_sc_hd__a211oi_4 _09843_ (.A1(_03242_),
    .A2(_03245_),
    .B1(_03480_),
    .C1(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__o211a_1 _09844_ (.A1(_03480_),
    .A2(_03481_),
    .B1(_03242_),
    .C1(_03245_),
    .X(_03483_));
 sky130_fd_sc_hd__a211oi_2 _09845_ (.A1(_03333_),
    .A2(_03335_),
    .B1(_03482_),
    .C1(_03483_),
    .Y(_03485_));
 sky130_fd_sc_hd__o211a_1 _09846_ (.A1(_03482_),
    .A2(_03483_),
    .B1(_03333_),
    .C1(_03335_),
    .X(_03486_));
 sky130_fd_sc_hd__a211oi_2 _09847_ (.A1(_03214_),
    .A2(_03217_),
    .B1(_03485_),
    .C1(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__o211a_1 _09848_ (.A1(_03485_),
    .A2(_03486_),
    .B1(_03214_),
    .C1(_03217_),
    .X(_03488_));
 sky130_fd_sc_hd__a211oi_1 _09849_ (.A1(_03337_),
    .A2(_03339_),
    .B1(_03487_),
    .C1(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__o211ai_2 _09850_ (.A1(_03487_),
    .A2(_03488_),
    .B1(_03337_),
    .C1(_03339_),
    .Y(_03490_));
 sky130_fd_sc_hd__nand2b_1 _09851_ (.A_N(_03489_),
    .B(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__a31o_1 _09852_ (.A1(_03339_),
    .A2(_03340_),
    .A3(_03342_),
    .B1(_03352_),
    .X(_03492_));
 sky130_fd_sc_hd__xnor2_1 _09853_ (.A(_03491_),
    .B(_03492_),
    .Y(net100));
 sky130_fd_sc_hd__nand2b_1 _09854_ (.A_N(_03390_),
    .B(_03392_),
    .Y(_03493_));
 sky130_fd_sc_hd__and4_1 _09855_ (.A(net6),
    .B(net7),
    .C(net52),
    .D(net53),
    .X(_03495_));
 sky130_fd_sc_hd__a22o_1 _09856_ (.A1(net7),
    .A2(net52),
    .B1(net53),
    .B2(net6),
    .X(_03496_));
 sky130_fd_sc_hd__and2b_1 _09857_ (.A_N(_03495_),
    .B(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__nand2_1 _09858_ (.A(net5),
    .B(net54),
    .Y(_03498_));
 sky130_fd_sc_hd__xnor2_1 _09859_ (.A(_03497_),
    .B(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__a31o_1 _09860_ (.A1(net4),
    .A2(net54),
    .A3(_03356_),
    .B1(_03355_),
    .X(_03500_));
 sky130_fd_sc_hd__nand2_1 _09861_ (.A(_03499_),
    .B(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__xor2_1 _09862_ (.A(_03499_),
    .B(_03500_),
    .X(_03502_));
 sky130_fd_sc_hd__and4b_1 _09863_ (.A_N(net3),
    .B(net4),
    .C(net56),
    .D(net57),
    .X(_03503_));
 sky130_fd_sc_hd__o2bb2a_1 _09864_ (.A1_N(net4),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net3),
    .X(_03504_));
 sky130_fd_sc_hd__nor2_1 _09865_ (.A(_03503_),
    .B(_03504_),
    .Y(_03506_));
 sky130_fd_sc_hd__xnor2_1 _09866_ (.A(_03502_),
    .B(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__a21bo_1 _09867_ (.A1(_03362_),
    .A2(_03365_),
    .B1_N(_03361_),
    .X(_03508_));
 sky130_fd_sc_hd__nand2b_1 _09868_ (.A_N(_03507_),
    .B(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__xor2_1 _09869_ (.A(_03507_),
    .B(_03508_),
    .X(_03510_));
 sky130_fd_sc_hd__inv_2 _09870_ (.A(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__nand2_1 _09871_ (.A(_03363_),
    .B(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__xor2_1 _09872_ (.A(_03363_),
    .B(_03510_),
    .X(_03513_));
 sky130_fd_sc_hd__a21o_1 _09873_ (.A1(_03404_),
    .A2(_03413_),
    .B1(_03412_),
    .X(_03514_));
 sky130_fd_sc_hd__nand2_1 _09874_ (.A(_03377_),
    .B(_03380_),
    .Y(_03515_));
 sky130_fd_sc_hd__a31o_1 _09875_ (.A1(net10),
    .A2(net48),
    .A3(_03401_),
    .B1(_03400_),
    .X(_03517_));
 sky130_fd_sc_hd__nand4_2 _09876_ (.A(net9),
    .B(net10),
    .C(net49),
    .D(net50),
    .Y(_03518_));
 sky130_fd_sc_hd__a22o_1 _09877_ (.A1(net10),
    .A2(net49),
    .B1(net50),
    .B2(net9),
    .X(_03519_));
 sky130_fd_sc_hd__a22o_1 _09878_ (.A1(net8),
    .A2(net51),
    .B1(_03518_),
    .B2(_03519_),
    .X(_03520_));
 sky130_fd_sc_hd__nand4_2 _09879_ (.A(net8),
    .B(net51),
    .C(_03518_),
    .D(_03519_),
    .Y(_03521_));
 sky130_fd_sc_hd__nand3_2 _09880_ (.A(_03517_),
    .B(_03520_),
    .C(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__a21o_1 _09881_ (.A1(_03520_),
    .A2(_03521_),
    .B1(_03517_),
    .X(_03523_));
 sky130_fd_sc_hd__nand3_2 _09882_ (.A(_03515_),
    .B(_03522_),
    .C(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__a21o_1 _09883_ (.A1(_03522_),
    .A2(_03523_),
    .B1(_03515_),
    .X(_03525_));
 sky130_fd_sc_hd__and3_1 _09884_ (.A(_03514_),
    .B(_03524_),
    .C(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__nand3_1 _09885_ (.A(_03514_),
    .B(_03524_),
    .C(_03525_),
    .Y(_03528_));
 sky130_fd_sc_hd__a21oi_1 _09886_ (.A1(_03524_),
    .A2(_03525_),
    .B1(_03514_),
    .Y(_03529_));
 sky130_fd_sc_hd__a211o_1 _09887_ (.A1(_03381_),
    .A2(_03383_),
    .B1(_03526_),
    .C1(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__o211ai_2 _09888_ (.A1(_03526_),
    .A2(_03529_),
    .B1(_03381_),
    .C1(_03383_),
    .Y(_03531_));
 sky130_fd_sc_hd__o211a_1 _09889_ (.A1(_03386_),
    .A2(_03388_),
    .B1(_03530_),
    .C1(_03531_),
    .X(_03532_));
 sky130_fd_sc_hd__a211oi_2 _09890_ (.A1(_03530_),
    .A2(_03531_),
    .B1(_03386_),
    .C1(_03388_),
    .Y(_03533_));
 sky130_fd_sc_hd__nor3_1 _09891_ (.A(_03513_),
    .B(_03532_),
    .C(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__or3_2 _09892_ (.A(_03513_),
    .B(_03532_),
    .C(_03533_),
    .X(_03535_));
 sky130_fd_sc_hd__o21ai_2 _09893_ (.A1(_03532_),
    .A2(_03533_),
    .B1(_03513_),
    .Y(_03536_));
 sky130_fd_sc_hd__o211ai_4 _09894_ (.A1(_03435_),
    .A2(_03437_),
    .B1(_03535_),
    .C1(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__a211o_1 _09895_ (.A1(_03535_),
    .A2(_03536_),
    .B1(_03435_),
    .C1(_03437_),
    .X(_03539_));
 sky130_fd_sc_hd__nand3_2 _09896_ (.A(_03493_),
    .B(_03537_),
    .C(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__a21o_1 _09897_ (.A1(_03537_),
    .A2(_03539_),
    .B1(_03493_),
    .X(_03541_));
 sky130_fd_sc_hd__and4_1 _09898_ (.A(net13),
    .B(net14),
    .C(net46),
    .D(net47),
    .X(_03542_));
 sky130_fd_sc_hd__a22o_1 _09899_ (.A1(net14),
    .A2(net46),
    .B1(net47),
    .B2(net13),
    .X(_03543_));
 sky130_fd_sc_hd__and2b_1 _09900_ (.A_N(_03542_),
    .B(_03543_),
    .X(_03544_));
 sky130_fd_sc_hd__nand2_1 _09901_ (.A(net11),
    .B(net48),
    .Y(_03545_));
 sky130_fd_sc_hd__xnor2_2 _09902_ (.A(_03544_),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__nand4_1 _09903_ (.A(net42),
    .B(net43),
    .C(net16),
    .D(net17),
    .Y(_03547_));
 sky130_fd_sc_hd__a22o_1 _09904_ (.A1(net43),
    .A2(net16),
    .B1(net17),
    .B2(net42),
    .X(_03548_));
 sky130_fd_sc_hd__and2_1 _09905_ (.A(net45),
    .B(net15),
    .X(_03550_));
 sky130_fd_sc_hd__a21o_1 _09906_ (.A1(_03547_),
    .A2(_03548_),
    .B1(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__nand3_1 _09907_ (.A(_03547_),
    .B(_03548_),
    .C(_03550_),
    .Y(_03552_));
 sky130_fd_sc_hd__a21bo_1 _09908_ (.A1(_03406_),
    .A2(_03408_),
    .B1_N(_03405_),
    .X(_03553_));
 sky130_fd_sc_hd__and3_1 _09909_ (.A(_03551_),
    .B(_03552_),
    .C(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__a21o_1 _09910_ (.A1(_03551_),
    .A2(_03552_),
    .B1(_03553_),
    .X(_03555_));
 sky130_fd_sc_hd__and2b_1 _09911_ (.A_N(_03554_),
    .B(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__xnor2_2 _09912_ (.A(_03546_),
    .B(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__nand2_1 _09913_ (.A(_03419_),
    .B(_03422_),
    .Y(_03558_));
 sky130_fd_sc_hd__a31o_1 _09914_ (.A1(net38),
    .A2(net20),
    .A3(_03444_),
    .B1(_03443_),
    .X(_03559_));
 sky130_fd_sc_hd__nand4_1 _09915_ (.A(net39),
    .B(net40),
    .C(net19),
    .D(net20),
    .Y(_03561_));
 sky130_fd_sc_hd__a22o_1 _09916_ (.A1(net40),
    .A2(net19),
    .B1(net20),
    .B2(net39),
    .X(_03562_));
 sky130_fd_sc_hd__a22o_1 _09917_ (.A1(net41),
    .A2(net18),
    .B1(_03561_),
    .B2(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__nand4_1 _09918_ (.A(net41),
    .B(net18),
    .C(_03561_),
    .D(_03562_),
    .Y(_03564_));
 sky130_fd_sc_hd__nand3_1 _09919_ (.A(_03559_),
    .B(_03563_),
    .C(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__a21o_1 _09920_ (.A1(_03563_),
    .A2(_03564_),
    .B1(_03559_),
    .X(_03566_));
 sky130_fd_sc_hd__nand3_1 _09921_ (.A(_03558_),
    .B(_03565_),
    .C(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__a21o_1 _09922_ (.A1(_03565_),
    .A2(_03566_),
    .B1(_03558_),
    .X(_03568_));
 sky130_fd_sc_hd__a21bo_1 _09923_ (.A1(_03416_),
    .A2(_03424_),
    .B1_N(_03423_),
    .X(_03569_));
 sky130_fd_sc_hd__and3_1 _09924_ (.A(_03567_),
    .B(_03568_),
    .C(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__a21oi_1 _09925_ (.A1(_03567_),
    .A2(_03568_),
    .B1(_03569_),
    .Y(_03572_));
 sky130_fd_sc_hd__nor3_2 _09926_ (.A(_03557_),
    .B(_03570_),
    .C(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__o21a_1 _09927_ (.A1(_03570_),
    .A2(_03572_),
    .B1(_03557_),
    .X(_03574_));
 sky130_fd_sc_hd__a211oi_4 _09928_ (.A1(_03458_),
    .A2(_03460_),
    .B1(_03573_),
    .C1(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__o211a_1 _09929_ (.A1(_03573_),
    .A2(_03574_),
    .B1(_03458_),
    .C1(_03460_),
    .X(_03576_));
 sky130_fd_sc_hd__a211oi_2 _09930_ (.A1(_03430_),
    .A2(_03433_),
    .B1(_03575_),
    .C1(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__o211a_1 _09931_ (.A1(_03575_),
    .A2(_03576_),
    .B1(_03430_),
    .C1(_03433_),
    .X(_03578_));
 sky130_fd_sc_hd__nand2_1 _09932_ (.A(_03454_),
    .B(_03456_),
    .Y(_03579_));
 sky130_fd_sc_hd__and4_1 _09933_ (.A(net36),
    .B(net37),
    .C(net22),
    .D(net24),
    .X(_03580_));
 sky130_fd_sc_hd__a22o_1 _09934_ (.A1(net37),
    .A2(net22),
    .B1(net24),
    .B2(net36),
    .X(_03581_));
 sky130_fd_sc_hd__and2b_1 _09935_ (.A_N(_03580_),
    .B(_03581_),
    .X(_03583_));
 sky130_fd_sc_hd__nand2_1 _09936_ (.A(net38),
    .B(net21),
    .Y(_03584_));
 sky130_fd_sc_hd__xnor2_1 _09937_ (.A(_03583_),
    .B(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__o21bai_1 _09938_ (.A1(_03448_),
    .A2(_03449_),
    .B1_N(_03294_),
    .Y(_03586_));
 sky130_fd_sc_hd__nand2_1 _09939_ (.A(net35),
    .B(net25),
    .Y(_03587_));
 sky130_fd_sc_hd__o21ai_1 _09940_ (.A1(_03294_),
    .A2(_03448_),
    .B1(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__or3_1 _09941_ (.A(_03294_),
    .B(_03448_),
    .C(_03587_),
    .X(_03589_));
 sky130_fd_sc_hd__and2_1 _09942_ (.A(net35),
    .B(_03294_),
    .X(_03590_));
 sky130_fd_sc_hd__nand2_2 _09943_ (.A(net35),
    .B(_03294_),
    .Y(_03591_));
 sky130_fd_sc_hd__a21o_1 _09944_ (.A1(_03588_),
    .A2(_03589_),
    .B1(_03586_),
    .X(_03592_));
 sky130_fd_sc_hd__and3_1 _09945_ (.A(_03585_),
    .B(_03591_),
    .C(_03592_),
    .X(_03594_));
 sky130_fd_sc_hd__a21oi_1 _09946_ (.A1(_03591_),
    .A2(_03592_),
    .B1(_03585_),
    .Y(_03595_));
 sky130_fd_sc_hd__or3_2 _09947_ (.A(_03441_),
    .B(_03594_),
    .C(_03595_),
    .X(_03596_));
 sky130_fd_sc_hd__o21ai_1 _09948_ (.A1(_03594_),
    .A2(_03595_),
    .B1(_03441_),
    .Y(_03597_));
 sky130_fd_sc_hd__nand3_2 _09949_ (.A(_03579_),
    .B(_03596_),
    .C(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__a21o_1 _09950_ (.A1(_03596_),
    .A2(_03597_),
    .B1(_03579_),
    .X(_03599_));
 sky130_fd_sc_hd__nand3_1 _09951_ (.A(_03465_),
    .B(_03598_),
    .C(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__a21o_1 _09952_ (.A1(_03598_),
    .A2(_03599_),
    .B1(_03465_),
    .X(_03601_));
 sky130_fd_sc_hd__a31o_1 _09953_ (.A1(_03460_),
    .A2(_03461_),
    .A3(_03465_),
    .B1(_03463_),
    .X(_03602_));
 sky130_fd_sc_hd__nand3_1 _09954_ (.A(_03600_),
    .B(_03601_),
    .C(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__a21o_1 _09955_ (.A1(_03600_),
    .A2(_03601_),
    .B1(_03602_),
    .X(_03605_));
 sky130_fd_sc_hd__or4bb_2 _09956_ (.A(_03577_),
    .B(_03578_),
    .C_N(_03603_),
    .D_N(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__a2bb2o_1 _09957_ (.A1_N(_03577_),
    .A2_N(_03578_),
    .B1(_03603_),
    .B2(_03605_),
    .X(_03607_));
 sky130_fd_sc_hd__o211ai_4 _09958_ (.A1(_03470_),
    .A2(_03472_),
    .B1(_03606_),
    .C1(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__inv_2 _09959_ (.A(_03608_),
    .Y(_03609_));
 sky130_fd_sc_hd__a211o_1 _09960_ (.A1(_03606_),
    .A2(_03607_),
    .B1(_03470_),
    .C1(_03472_),
    .X(_03610_));
 sky130_fd_sc_hd__and4_1 _09961_ (.A(_03540_),
    .B(_03541_),
    .C(_03608_),
    .D(_03610_),
    .X(_03611_));
 sky130_fd_sc_hd__nand4_2 _09962_ (.A(_03540_),
    .B(_03541_),
    .C(_03608_),
    .D(_03610_),
    .Y(_03612_));
 sky130_fd_sc_hd__a22o_1 _09963_ (.A1(_03540_),
    .A2(_03541_),
    .B1(_03608_),
    .B2(_03610_),
    .X(_03613_));
 sky130_fd_sc_hd__o211ai_4 _09964_ (.A1(_03476_),
    .A2(_03478_),
    .B1(_03612_),
    .C1(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__a211o_1 _09965_ (.A1(_03612_),
    .A2(_03613_),
    .B1(_03476_),
    .C1(_03478_),
    .X(_03616_));
 sky130_fd_sc_hd__o211ai_4 _09966_ (.A1(_03394_),
    .A2(_03398_),
    .B1(_03614_),
    .C1(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__a211o_1 _09967_ (.A1(_03614_),
    .A2(_03616_),
    .B1(_03394_),
    .C1(_03398_),
    .X(_03618_));
 sky130_fd_sc_hd__o211ai_4 _09968_ (.A1(_03480_),
    .A2(_03482_),
    .B1(_03617_),
    .C1(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__a211o_1 _09969_ (.A1(_03617_),
    .A2(_03618_),
    .B1(_03480_),
    .C1(_03482_),
    .X(_03620_));
 sky130_fd_sc_hd__o211ai_2 _09970_ (.A1(_03368_),
    .A2(_03371_),
    .B1(_03619_),
    .C1(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__a211o_1 _09971_ (.A1(_03619_),
    .A2(_03620_),
    .B1(_03368_),
    .C1(_03371_),
    .X(_03622_));
 sky130_fd_sc_hd__o211a_1 _09972_ (.A1(_03485_),
    .A2(_03487_),
    .B1(_03621_),
    .C1(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__a211oi_1 _09973_ (.A1(_03621_),
    .A2(_03622_),
    .B1(_03485_),
    .C1(_03487_),
    .Y(_03624_));
 sky130_fd_sc_hd__nor2_1 _09974_ (.A(_03623_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__a41oi_2 _09975_ (.A1(_03339_),
    .A2(_03340_),
    .A3(_03342_),
    .A4(_03490_),
    .B1(_03489_),
    .Y(_03627_));
 sky130_fd_sc_hd__o31a_1 _09976_ (.A1(_03344_),
    .A2(_03351_),
    .A3(_03491_),
    .B1(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__xnor2_1 _09977_ (.A(_03625_),
    .B(_03628_),
    .Y(net101));
 sky130_fd_sc_hd__and4_1 _09978_ (.A(net7),
    .B(net8),
    .C(net52),
    .D(net53),
    .X(_03629_));
 sky130_fd_sc_hd__a22o_1 _09979_ (.A1(net8),
    .A2(net52),
    .B1(net53),
    .B2(net7),
    .X(_03630_));
 sky130_fd_sc_hd__and2b_1 _09980_ (.A_N(_03629_),
    .B(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__nand2_1 _09981_ (.A(net6),
    .B(net54),
    .Y(_03632_));
 sky130_fd_sc_hd__xnor2_1 _09982_ (.A(_03631_),
    .B(_03632_),
    .Y(_03633_));
 sky130_fd_sc_hd__a31o_1 _09983_ (.A1(net5),
    .A2(net54),
    .A3(_03496_),
    .B1(_03495_),
    .X(_03634_));
 sky130_fd_sc_hd__nand2_1 _09984_ (.A(_03633_),
    .B(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__xor2_1 _09985_ (.A(_03633_),
    .B(_03634_),
    .X(_03637_));
 sky130_fd_sc_hd__and4b_1 _09986_ (.A_N(net4),
    .B(net5),
    .C(net56),
    .D(net57),
    .X(_03638_));
 sky130_fd_sc_hd__o2bb2a_1 _09987_ (.A1_N(net5),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net4),
    .X(_03639_));
 sky130_fd_sc_hd__nor2_1 _09988_ (.A(_03638_),
    .B(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__xnor2_1 _09989_ (.A(_03637_),
    .B(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__a21bo_1 _09990_ (.A1(_03502_),
    .A2(_03506_),
    .B1_N(_03501_),
    .X(_03642_));
 sky130_fd_sc_hd__and2b_1 _09991_ (.A_N(_03641_),
    .B(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__xor2_1 _09992_ (.A(_03641_),
    .B(_03642_),
    .X(_03644_));
 sky130_fd_sc_hd__inv_2 _09993_ (.A(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__xor2_1 _09994_ (.A(_03503_),
    .B(_03644_),
    .X(_03646_));
 sky130_fd_sc_hd__a21o_1 _09995_ (.A1(_03546_),
    .A2(_03555_),
    .B1(_03554_),
    .X(_03648_));
 sky130_fd_sc_hd__nand2_1 _09996_ (.A(_03518_),
    .B(_03521_),
    .Y(_03649_));
 sky130_fd_sc_hd__a31o_1 _09997_ (.A1(net11),
    .A2(net48),
    .A3(_03543_),
    .B1(_03542_),
    .X(_03650_));
 sky130_fd_sc_hd__nand4_2 _09998_ (.A(net10),
    .B(net11),
    .C(net49),
    .D(net50),
    .Y(_03651_));
 sky130_fd_sc_hd__a22o_1 _09999_ (.A1(net11),
    .A2(net49),
    .B1(net50),
    .B2(net10),
    .X(_03652_));
 sky130_fd_sc_hd__a22o_1 _10000_ (.A1(net9),
    .A2(net51),
    .B1(_03651_),
    .B2(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__nand4_2 _10001_ (.A(net9),
    .B(net51),
    .C(_03651_),
    .D(_03652_),
    .Y(_03654_));
 sky130_fd_sc_hd__nand3_2 _10002_ (.A(_03650_),
    .B(_03653_),
    .C(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__a21o_1 _10003_ (.A1(_03653_),
    .A2(_03654_),
    .B1(_03650_),
    .X(_03656_));
 sky130_fd_sc_hd__nand3_2 _10004_ (.A(_03649_),
    .B(_03655_),
    .C(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__a21o_1 _10005_ (.A1(_03655_),
    .A2(_03656_),
    .B1(_03649_),
    .X(_03659_));
 sky130_fd_sc_hd__and3_1 _10006_ (.A(_03648_),
    .B(_03657_),
    .C(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__a21oi_1 _10007_ (.A1(_03657_),
    .A2(_03659_),
    .B1(_03648_),
    .Y(_03661_));
 sky130_fd_sc_hd__a211oi_2 _10008_ (.A1(_03522_),
    .A2(_03524_),
    .B1(_03660_),
    .C1(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__o211a_1 _10009_ (.A1(_03660_),
    .A2(_03661_),
    .B1(_03522_),
    .C1(_03524_),
    .X(_03663_));
 sky130_fd_sc_hd__a211oi_1 _10010_ (.A1(_03528_),
    .A2(_03530_),
    .B1(_03662_),
    .C1(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__o211a_1 _10011_ (.A1(_03662_),
    .A2(_03663_),
    .B1(_03528_),
    .C1(_03530_),
    .X(_03665_));
 sky130_fd_sc_hd__or3_1 _10012_ (.A(_03646_),
    .B(_03664_),
    .C(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__o21ai_1 _10013_ (.A1(_03664_),
    .A2(_03665_),
    .B1(_03646_),
    .Y(_03667_));
 sky130_fd_sc_hd__o211a_1 _10014_ (.A1(_03575_),
    .A2(_03577_),
    .B1(_03666_),
    .C1(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__o211ai_1 _10015_ (.A1(_03575_),
    .A2(_03577_),
    .B1(_03666_),
    .C1(_03667_),
    .Y(_03670_));
 sky130_fd_sc_hd__a211o_1 _10016_ (.A1(_03666_),
    .A2(_03667_),
    .B1(_03575_),
    .C1(_03577_),
    .X(_03671_));
 sky130_fd_sc_hd__o211a_1 _10017_ (.A1(_03532_),
    .A2(_03534_),
    .B1(_03670_),
    .C1(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__a211oi_1 _10018_ (.A1(_03670_),
    .A2(_03671_),
    .B1(_03532_),
    .C1(_03534_),
    .Y(_03673_));
 sky130_fd_sc_hd__and4_1 _10019_ (.A(net14),
    .B(net46),
    .C(net15),
    .D(net47),
    .X(_03674_));
 sky130_fd_sc_hd__a22o_1 _10020_ (.A1(net46),
    .A2(net15),
    .B1(net47),
    .B2(net14),
    .X(_03675_));
 sky130_fd_sc_hd__and2b_1 _10021_ (.A_N(_03674_),
    .B(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__nand2_1 _10022_ (.A(net13),
    .B(net48),
    .Y(_03677_));
 sky130_fd_sc_hd__xnor2_2 _10023_ (.A(_03676_),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__nand4_1 _10024_ (.A(net42),
    .B(net43),
    .C(net17),
    .D(net18),
    .Y(_03679_));
 sky130_fd_sc_hd__a22o_1 _10025_ (.A1(net43),
    .A2(net17),
    .B1(net18),
    .B2(net42),
    .X(_03681_));
 sky130_fd_sc_hd__and2_1 _10026_ (.A(net45),
    .B(net16),
    .X(_03682_));
 sky130_fd_sc_hd__a21o_1 _10027_ (.A1(_03679_),
    .A2(_03681_),
    .B1(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__nand3_1 _10028_ (.A(_03679_),
    .B(_03681_),
    .C(_03682_),
    .Y(_03684_));
 sky130_fd_sc_hd__a21bo_1 _10029_ (.A1(_03548_),
    .A2(_03550_),
    .B1_N(_03547_),
    .X(_03685_));
 sky130_fd_sc_hd__and3_1 _10030_ (.A(_03683_),
    .B(_03684_),
    .C(_03685_),
    .X(_03686_));
 sky130_fd_sc_hd__a21o_1 _10031_ (.A1(_03683_),
    .A2(_03684_),
    .B1(_03685_),
    .X(_03687_));
 sky130_fd_sc_hd__and2b_1 _10032_ (.A_N(_03686_),
    .B(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__xnor2_2 _10033_ (.A(_03678_),
    .B(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__nand2_1 _10034_ (.A(_03561_),
    .B(_03564_),
    .Y(_03690_));
 sky130_fd_sc_hd__a31o_1 _10035_ (.A1(net38),
    .A2(net21),
    .A3(_03581_),
    .B1(_03580_),
    .X(_03692_));
 sky130_fd_sc_hd__nand4_1 _10036_ (.A(net39),
    .B(net40),
    .C(net20),
    .D(net21),
    .Y(_03693_));
 sky130_fd_sc_hd__a22o_1 _10037_ (.A1(net40),
    .A2(net20),
    .B1(net21),
    .B2(net39),
    .X(_03694_));
 sky130_fd_sc_hd__a22o_1 _10038_ (.A1(net41),
    .A2(net19),
    .B1(_03693_),
    .B2(_03694_),
    .X(_03695_));
 sky130_fd_sc_hd__nand4_1 _10039_ (.A(net41),
    .B(net19),
    .C(_03693_),
    .D(_03694_),
    .Y(_03696_));
 sky130_fd_sc_hd__nand3_1 _10040_ (.A(_03692_),
    .B(_03695_),
    .C(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__a21o_1 _10041_ (.A1(_03695_),
    .A2(_03696_),
    .B1(_03692_),
    .X(_03698_));
 sky130_fd_sc_hd__nand3_1 _10042_ (.A(_03690_),
    .B(_03697_),
    .C(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__a21o_1 _10043_ (.A1(_03697_),
    .A2(_03698_),
    .B1(_03690_),
    .X(_03700_));
 sky130_fd_sc_hd__a21bo_1 _10044_ (.A1(_03558_),
    .A2(_03566_),
    .B1_N(_03565_),
    .X(_03701_));
 sky130_fd_sc_hd__and3_2 _10045_ (.A(_03699_),
    .B(_03700_),
    .C(_03701_),
    .X(_03703_));
 sky130_fd_sc_hd__a21oi_1 _10046_ (.A1(_03699_),
    .A2(_03700_),
    .B1(_03701_),
    .Y(_03704_));
 sky130_fd_sc_hd__nor3_2 _10047_ (.A(_03689_),
    .B(_03703_),
    .C(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__o21a_1 _10048_ (.A1(_03703_),
    .A2(_03704_),
    .B1(_03689_),
    .X(_03706_));
 sky130_fd_sc_hd__a211o_1 _10049_ (.A1(_03596_),
    .A2(_03598_),
    .B1(_03705_),
    .C1(_03706_),
    .X(_03707_));
 sky130_fd_sc_hd__o211ai_2 _10050_ (.A1(_03705_),
    .A2(_03706_),
    .B1(_03596_),
    .C1(_03598_),
    .Y(_03708_));
 sky130_fd_sc_hd__o211ai_2 _10051_ (.A1(_03570_),
    .A2(_03573_),
    .B1(_03707_),
    .C1(_03708_),
    .Y(_03709_));
 sky130_fd_sc_hd__a211o_1 _10052_ (.A1(_03707_),
    .A2(_03708_),
    .B1(_03570_),
    .C1(_03573_),
    .X(_03710_));
 sky130_fd_sc_hd__nor2_1 _10053_ (.A(_03590_),
    .B(_03594_),
    .Y(_03711_));
 sky130_fd_sc_hd__and4_1 _10054_ (.A(net36),
    .B(net37),
    .C(net24),
    .D(net25),
    .X(_03712_));
 sky130_fd_sc_hd__a22o_1 _10055_ (.A1(net37),
    .A2(net24),
    .B1(net25),
    .B2(net36),
    .X(_03714_));
 sky130_fd_sc_hd__nand2b_1 _10056_ (.A_N(_03712_),
    .B(_03714_),
    .Y(_03715_));
 sky130_fd_sc_hd__nand2_1 _10057_ (.A(net38),
    .B(net22),
    .Y(_03716_));
 sky130_fd_sc_hd__xnor2_1 _10058_ (.A(_03715_),
    .B(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__a21o_2 _10059_ (.A1(_03448_),
    .A2(_03587_),
    .B1(_03590_),
    .X(_03718_));
 sky130_fd_sc_hd__xnor2_1 _10060_ (.A(_03717_),
    .B(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__nor2_1 _10061_ (.A(_03441_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__xnor2_1 _10062_ (.A(_03442_),
    .B(_03719_),
    .Y(_03721_));
 sky130_fd_sc_hd__and2b_1 _10063_ (.A_N(_03711_),
    .B(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__xnor2_1 _10064_ (.A(_03711_),
    .B(_03721_),
    .Y(_03723_));
 sky130_fd_sc_hd__xnor2_1 _10065_ (.A(_03465_),
    .B(_03723_),
    .Y(_03725_));
 sky130_fd_sc_hd__a31o_1 _10066_ (.A1(_03465_),
    .A2(_03598_),
    .A3(_03599_),
    .B1(_03463_),
    .X(_03726_));
 sky130_fd_sc_hd__and2b_1 _10067_ (.A_N(_03725_),
    .B(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__xnor2_1 _10068_ (.A(_03725_),
    .B(_03726_),
    .Y(_03728_));
 sky130_fd_sc_hd__and3_1 _10069_ (.A(_03709_),
    .B(_03710_),
    .C(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__a21oi_1 _10070_ (.A1(_03709_),
    .A2(_03710_),
    .B1(_03728_),
    .Y(_03730_));
 sky130_fd_sc_hd__a211o_1 _10071_ (.A1(_03603_),
    .A2(_03606_),
    .B1(_03729_),
    .C1(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__o211ai_1 _10072_ (.A1(_03729_),
    .A2(_03730_),
    .B1(_03603_),
    .C1(_03606_),
    .Y(_03732_));
 sky130_fd_sc_hd__or4bb_2 _10073_ (.A(_03672_),
    .B(_03673_),
    .C_N(_03731_),
    .D_N(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__a2bb2o_1 _10074_ (.A1_N(_03672_),
    .A2_N(_03673_),
    .B1(_03731_),
    .B2(_03732_),
    .X(_03734_));
 sky130_fd_sc_hd__o211a_1 _10075_ (.A1(_03609_),
    .A2(_03611_),
    .B1(_03733_),
    .C1(_03734_),
    .X(_03736_));
 sky130_fd_sc_hd__a211oi_1 _10076_ (.A1(_03733_),
    .A2(_03734_),
    .B1(_03609_),
    .C1(_03611_),
    .Y(_03737_));
 sky130_fd_sc_hd__a211oi_2 _10077_ (.A1(_03537_),
    .A2(_03540_),
    .B1(_03736_),
    .C1(_03737_),
    .Y(_03738_));
 sky130_fd_sc_hd__o211a_1 _10078_ (.A1(_03736_),
    .A2(_03737_),
    .B1(_03537_),
    .C1(_03540_),
    .X(_03739_));
 sky130_fd_sc_hd__a211oi_1 _10079_ (.A1(_03614_),
    .A2(_03617_),
    .B1(_03738_),
    .C1(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__o211a_1 _10080_ (.A1(_03738_),
    .A2(_03739_),
    .B1(_03614_),
    .C1(_03617_),
    .X(_03741_));
 sky130_fd_sc_hd__a211oi_1 _10081_ (.A1(_03509_),
    .A2(_03512_),
    .B1(_03740_),
    .C1(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__o211a_1 _10082_ (.A1(_03740_),
    .A2(_03741_),
    .B1(_03509_),
    .C1(_03512_),
    .X(_03743_));
 sky130_fd_sc_hd__o211ai_1 _10083_ (.A1(_03742_),
    .A2(_03743_),
    .B1(_03619_),
    .C1(_03621_),
    .Y(_03744_));
 sky130_fd_sc_hd__a211o_1 _10084_ (.A1(_03619_),
    .A2(_03621_),
    .B1(_03742_),
    .C1(_03743_),
    .X(_03745_));
 sky130_fd_sc_hd__and2_1 _10085_ (.A(_03744_),
    .B(_03745_),
    .X(_03747_));
 sky130_fd_sc_hd__o21ba_1 _10086_ (.A1(_03624_),
    .A2(_03628_),
    .B1_N(_03623_),
    .X(_03748_));
 sky130_fd_sc_hd__xnor2_1 _10087_ (.A(_03747_),
    .B(_03748_),
    .Y(net102));
 sky130_fd_sc_hd__a21oi_2 _10088_ (.A1(_03503_),
    .A2(_03645_),
    .B1(_03643_),
    .Y(_03749_));
 sky130_fd_sc_hd__nand2b_1 _10089_ (.A_N(_03664_),
    .B(_03666_),
    .Y(_03750_));
 sky130_fd_sc_hd__and4_1 _10090_ (.A(net8),
    .B(net9),
    .C(net52),
    .D(net53),
    .X(_03751_));
 sky130_fd_sc_hd__a22o_1 _10091_ (.A1(net9),
    .A2(net52),
    .B1(net53),
    .B2(net8),
    .X(_03752_));
 sky130_fd_sc_hd__and2b_1 _10092_ (.A_N(_03751_),
    .B(_03752_),
    .X(_03753_));
 sky130_fd_sc_hd__nand2_1 _10093_ (.A(net7),
    .B(net54),
    .Y(_03754_));
 sky130_fd_sc_hd__xnor2_1 _10094_ (.A(_03753_),
    .B(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__a31o_1 _10095_ (.A1(net6),
    .A2(net54),
    .A3(_03630_),
    .B1(_03629_),
    .X(_03757_));
 sky130_fd_sc_hd__nand2_1 _10096_ (.A(_03755_),
    .B(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__xor2_1 _10097_ (.A(_03755_),
    .B(_03757_),
    .X(_03759_));
 sky130_fd_sc_hd__and4b_1 _10098_ (.A_N(net5),
    .B(net6),
    .C(net56),
    .D(net57),
    .X(_03760_));
 sky130_fd_sc_hd__o2bb2a_1 _10099_ (.A1_N(net6),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net5),
    .X(_03761_));
 sky130_fd_sc_hd__nor2_1 _10100_ (.A(_03760_),
    .B(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__xnor2_1 _10101_ (.A(_03759_),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__a21bo_1 _10102_ (.A1(_03637_),
    .A2(_03640_),
    .B1_N(_03635_),
    .X(_03764_));
 sky130_fd_sc_hd__nand2b_1 _10103_ (.A_N(_03763_),
    .B(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__xor2_1 _10104_ (.A(_03763_),
    .B(_03764_),
    .X(_03766_));
 sky130_fd_sc_hd__inv_2 _10105_ (.A(_03766_),
    .Y(_03768_));
 sky130_fd_sc_hd__nand2_1 _10106_ (.A(_03638_),
    .B(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__xor2_1 _10107_ (.A(_03638_),
    .B(_03766_),
    .X(_03770_));
 sky130_fd_sc_hd__a21o_1 _10108_ (.A1(_03678_),
    .A2(_03687_),
    .B1(_03686_),
    .X(_03771_));
 sky130_fd_sc_hd__nand2_1 _10109_ (.A(_03651_),
    .B(_03654_),
    .Y(_03772_));
 sky130_fd_sc_hd__a31o_1 _10110_ (.A1(net13),
    .A2(net48),
    .A3(_03675_),
    .B1(_03674_),
    .X(_03773_));
 sky130_fd_sc_hd__nand4_2 _10111_ (.A(net11),
    .B(net13),
    .C(net49),
    .D(net50),
    .Y(_03774_));
 sky130_fd_sc_hd__a22o_1 _10112_ (.A1(net13),
    .A2(net49),
    .B1(net50),
    .B2(net11),
    .X(_03775_));
 sky130_fd_sc_hd__a22o_1 _10113_ (.A1(net10),
    .A2(net51),
    .B1(_03774_),
    .B2(_03775_),
    .X(_03776_));
 sky130_fd_sc_hd__nand4_2 _10114_ (.A(net10),
    .B(net51),
    .C(_03774_),
    .D(_03775_),
    .Y(_03777_));
 sky130_fd_sc_hd__nand3_2 _10115_ (.A(_03773_),
    .B(_03776_),
    .C(_03777_),
    .Y(_03779_));
 sky130_fd_sc_hd__a21o_1 _10116_ (.A1(_03776_),
    .A2(_03777_),
    .B1(_03773_),
    .X(_03780_));
 sky130_fd_sc_hd__nand3_2 _10117_ (.A(_03772_),
    .B(_03779_),
    .C(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__a21o_1 _10118_ (.A1(_03779_),
    .A2(_03780_),
    .B1(_03772_),
    .X(_03782_));
 sky130_fd_sc_hd__and3_1 _10119_ (.A(_03771_),
    .B(_03781_),
    .C(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__nand3_1 _10120_ (.A(_03771_),
    .B(_03781_),
    .C(_03782_),
    .Y(_03784_));
 sky130_fd_sc_hd__a21oi_1 _10121_ (.A1(_03781_),
    .A2(_03782_),
    .B1(_03771_),
    .Y(_03785_));
 sky130_fd_sc_hd__a211o_1 _10122_ (.A1(_03655_),
    .A2(_03657_),
    .B1(_03783_),
    .C1(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__o211ai_2 _10123_ (.A1(_03783_),
    .A2(_03785_),
    .B1(_03655_),
    .C1(_03657_),
    .Y(_03787_));
 sky130_fd_sc_hd__o211a_1 _10124_ (.A1(_03660_),
    .A2(_03662_),
    .B1(_03786_),
    .C1(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__a211oi_2 _10125_ (.A1(_03786_),
    .A2(_03787_),
    .B1(_03660_),
    .C1(_03662_),
    .Y(_03790_));
 sky130_fd_sc_hd__nor3_2 _10126_ (.A(_03770_),
    .B(_03788_),
    .C(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__o21a_1 _10127_ (.A1(_03788_),
    .A2(_03790_),
    .B1(_03770_),
    .X(_03792_));
 sky130_fd_sc_hd__a211o_2 _10128_ (.A1(_03707_),
    .A2(_03709_),
    .B1(_03791_),
    .C1(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__o211ai_2 _10129_ (.A1(_03791_),
    .A2(_03792_),
    .B1(_03707_),
    .C1(_03709_),
    .Y(_03794_));
 sky130_fd_sc_hd__nand3_2 _10130_ (.A(_03750_),
    .B(_03793_),
    .C(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__a21o_1 _10131_ (.A1(_03793_),
    .A2(_03794_),
    .B1(_03750_),
    .X(_03796_));
 sky130_fd_sc_hd__and4_1 _10132_ (.A(net46),
    .B(net15),
    .C(net47),
    .D(net16),
    .X(_03797_));
 sky130_fd_sc_hd__a22o_1 _10133_ (.A1(net15),
    .A2(net47),
    .B1(net16),
    .B2(net46),
    .X(_03798_));
 sky130_fd_sc_hd__and2b_1 _10134_ (.A_N(_03797_),
    .B(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__nand2_1 _10135_ (.A(net14),
    .B(net48),
    .Y(_03801_));
 sky130_fd_sc_hd__xnor2_1 _10136_ (.A(_03799_),
    .B(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__nand4_1 _10137_ (.A(net42),
    .B(net43),
    .C(net18),
    .D(net19),
    .Y(_03803_));
 sky130_fd_sc_hd__a22o_1 _10138_ (.A1(net43),
    .A2(net18),
    .B1(net19),
    .B2(net42),
    .X(_03804_));
 sky130_fd_sc_hd__and2_1 _10139_ (.A(net45),
    .B(net17),
    .X(_03805_));
 sky130_fd_sc_hd__a21o_1 _10140_ (.A1(_03803_),
    .A2(_03804_),
    .B1(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__nand3_1 _10141_ (.A(_03803_),
    .B(_03804_),
    .C(_03805_),
    .Y(_03807_));
 sky130_fd_sc_hd__a21bo_1 _10142_ (.A1(_03681_),
    .A2(_03682_),
    .B1_N(_03679_),
    .X(_03808_));
 sky130_fd_sc_hd__and3_1 _10143_ (.A(_03806_),
    .B(_03807_),
    .C(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__a21o_1 _10144_ (.A1(_03806_),
    .A2(_03807_),
    .B1(_03808_),
    .X(_03810_));
 sky130_fd_sc_hd__and2b_1 _10145_ (.A_N(_03809_),
    .B(_03810_),
    .X(_03812_));
 sky130_fd_sc_hd__xnor2_1 _10146_ (.A(_03802_),
    .B(_03812_),
    .Y(_03813_));
 sky130_fd_sc_hd__nand2_1 _10147_ (.A(_03693_),
    .B(_03696_),
    .Y(_03814_));
 sky130_fd_sc_hd__a31o_1 _10148_ (.A1(net38),
    .A2(net22),
    .A3(_03714_),
    .B1(_03712_),
    .X(_03815_));
 sky130_fd_sc_hd__nand4_1 _10149_ (.A(net39),
    .B(net40),
    .C(net21),
    .D(net22),
    .Y(_03816_));
 sky130_fd_sc_hd__a22o_1 _10150_ (.A1(net40),
    .A2(net21),
    .B1(net22),
    .B2(net39),
    .X(_03817_));
 sky130_fd_sc_hd__a22o_1 _10151_ (.A1(net41),
    .A2(net20),
    .B1(_03816_),
    .B2(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__nand4_1 _10152_ (.A(net41),
    .B(net20),
    .C(_03816_),
    .D(_03817_),
    .Y(_03819_));
 sky130_fd_sc_hd__nand3_1 _10153_ (.A(_03815_),
    .B(_03818_),
    .C(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__a21o_1 _10154_ (.A1(_03818_),
    .A2(_03819_),
    .B1(_03815_),
    .X(_03821_));
 sky130_fd_sc_hd__nand3_1 _10155_ (.A(_03814_),
    .B(_03820_),
    .C(_03821_),
    .Y(_03823_));
 sky130_fd_sc_hd__a21o_1 _10156_ (.A1(_03820_),
    .A2(_03821_),
    .B1(_03814_),
    .X(_03824_));
 sky130_fd_sc_hd__a21bo_1 _10157_ (.A1(_03690_),
    .A2(_03698_),
    .B1_N(_03697_),
    .X(_03825_));
 sky130_fd_sc_hd__and3_1 _10158_ (.A(_03823_),
    .B(_03824_),
    .C(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__a21oi_1 _10159_ (.A1(_03823_),
    .A2(_03824_),
    .B1(_03825_),
    .Y(_03827_));
 sky130_fd_sc_hd__or3_2 _10160_ (.A(_03813_),
    .B(_03826_),
    .C(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__inv_2 _10161_ (.A(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__o21ai_2 _10162_ (.A1(_03826_),
    .A2(_03827_),
    .B1(_03813_),
    .Y(_03830_));
 sky130_fd_sc_hd__o211ai_4 _10163_ (.A1(_03720_),
    .A2(_03722_),
    .B1(_03828_),
    .C1(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__a211o_1 _10164_ (.A1(_03828_),
    .A2(_03830_),
    .B1(_03720_),
    .C1(_03722_),
    .X(_03832_));
 sky130_fd_sc_hd__o211ai_4 _10165_ (.A1(_03703_),
    .A2(_03705_),
    .B1(_03831_),
    .C1(_03832_),
    .Y(_03834_));
 sky130_fd_sc_hd__a211o_1 _10166_ (.A1(_03831_),
    .A2(_03832_),
    .B1(_03703_),
    .C1(_03705_),
    .X(_03835_));
 sky130_fd_sc_hd__o21ai_1 _10167_ (.A1(_03717_),
    .A2(_03718_),
    .B1(_03591_),
    .Y(_03836_));
 sky130_fd_sc_hd__and3_1 _10168_ (.A(net36),
    .B(net37),
    .C(net25),
    .X(_03837_));
 sky130_fd_sc_hd__o21a_1 _10169_ (.A1(net36),
    .A2(net37),
    .B1(net25),
    .X(_03838_));
 sky130_fd_sc_hd__and2b_2 _10170_ (.A_N(_03837_),
    .B(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__nand2_1 _10171_ (.A(net38),
    .B(net24),
    .Y(_03840_));
 sky130_fd_sc_hd__xor2_1 _10172_ (.A(_03839_),
    .B(_03840_),
    .X(_03841_));
 sky130_fd_sc_hd__xor2_1 _10173_ (.A(_03718_),
    .B(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__and2_1 _10174_ (.A(_03442_),
    .B(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__xnor2_1 _10175_ (.A(_03441_),
    .B(_03842_),
    .Y(_03845_));
 sky130_fd_sc_hd__and2_1 _10176_ (.A(_03836_),
    .B(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__xnor2_1 _10177_ (.A(_03836_),
    .B(_03845_),
    .Y(_03847_));
 sky130_fd_sc_hd__xnor2_1 _10178_ (.A(_03465_),
    .B(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__a21o_1 _10179_ (.A1(_03465_),
    .A2(_03723_),
    .B1(_03463_),
    .X(_03849_));
 sky130_fd_sc_hd__nand2_1 _10180_ (.A(_03848_),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__xor2_1 _10181_ (.A(_03848_),
    .B(_03849_),
    .X(_03851_));
 sky130_fd_sc_hd__nand3_2 _10182_ (.A(_03834_),
    .B(_03835_),
    .C(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__a21o_1 _10183_ (.A1(_03834_),
    .A2(_03835_),
    .B1(_03851_),
    .X(_03853_));
 sky130_fd_sc_hd__o211a_1 _10184_ (.A1(_03727_),
    .A2(_03729_),
    .B1(_03852_),
    .C1(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__o211ai_1 _10185_ (.A1(_03727_),
    .A2(_03729_),
    .B1(_03852_),
    .C1(_03853_),
    .Y(_03856_));
 sky130_fd_sc_hd__a211o_1 _10186_ (.A1(_03852_),
    .A2(_03853_),
    .B1(_03727_),
    .C1(_03729_),
    .X(_03857_));
 sky130_fd_sc_hd__and4_1 _10187_ (.A(_03795_),
    .B(_03796_),
    .C(_03856_),
    .D(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__a22oi_2 _10188_ (.A1(_03795_),
    .A2(_03796_),
    .B1(_03856_),
    .B2(_03857_),
    .Y(_03859_));
 sky130_fd_sc_hd__a211o_2 _10189_ (.A1(_03731_),
    .A2(_03733_),
    .B1(_03858_),
    .C1(_03859_),
    .X(_03860_));
 sky130_fd_sc_hd__o211ai_2 _10190_ (.A1(_03858_),
    .A2(_03859_),
    .B1(_03731_),
    .C1(_03733_),
    .Y(_03861_));
 sky130_fd_sc_hd__o211ai_4 _10191_ (.A1(_03668_),
    .A2(_03672_),
    .B1(_03860_),
    .C1(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__a211o_1 _10192_ (.A1(_03860_),
    .A2(_03861_),
    .B1(_03668_),
    .C1(_03672_),
    .X(_03863_));
 sky130_fd_sc_hd__o211a_1 _10193_ (.A1(_03736_),
    .A2(_03738_),
    .B1(_03862_),
    .C1(_03863_),
    .X(_03864_));
 sky130_fd_sc_hd__a211oi_1 _10194_ (.A1(_03862_),
    .A2(_03863_),
    .B1(_03736_),
    .C1(_03738_),
    .Y(_03865_));
 sky130_fd_sc_hd__or2_1 _10195_ (.A(_03864_),
    .B(_03865_),
    .X(_03867_));
 sky130_fd_sc_hd__xnor2_2 _10196_ (.A(_03749_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__nor2_1 _10197_ (.A(_03740_),
    .B(_03742_),
    .Y(_03869_));
 sky130_fd_sc_hd__xnor2_1 _10198_ (.A(_03868_),
    .B(_03869_),
    .Y(_03870_));
 sky130_fd_sc_hd__nand2_1 _10199_ (.A(_03625_),
    .B(_03747_),
    .Y(_03871_));
 sky130_fd_sc_hd__nand2_1 _10200_ (.A(_03623_),
    .B(_03744_),
    .Y(_03872_));
 sky130_fd_sc_hd__o211a_1 _10201_ (.A1(_03627_),
    .A2(_03871_),
    .B1(_03872_),
    .C1(_03745_),
    .X(_03873_));
 sky130_fd_sc_hd__nor2_1 _10202_ (.A(_03491_),
    .B(_03871_),
    .Y(_03874_));
 sky130_fd_sc_hd__a21boi_1 _10203_ (.A1(_03352_),
    .A2(_03874_),
    .B1_N(_03873_),
    .Y(_03875_));
 sky130_fd_sc_hd__or2_1 _10204_ (.A(_03870_),
    .B(_03875_),
    .X(_03876_));
 sky130_fd_sc_hd__nand2_1 _10205_ (.A(_03870_),
    .B(_03875_),
    .Y(_03878_));
 sky130_fd_sc_hd__and2_1 _10206_ (.A(_03876_),
    .B(_03878_),
    .X(net103));
 sky130_fd_sc_hd__o21ba_1 _10207_ (.A1(_03749_),
    .A2(_03865_),
    .B1_N(_03864_),
    .X(_03879_));
 sky130_fd_sc_hd__and4_1 _10208_ (.A(net9),
    .B(net10),
    .C(net52),
    .D(net53),
    .X(_03880_));
 sky130_fd_sc_hd__a22o_1 _10209_ (.A1(net10),
    .A2(net52),
    .B1(net53),
    .B2(net9),
    .X(_03881_));
 sky130_fd_sc_hd__and2b_1 _10210_ (.A_N(_03880_),
    .B(_03881_),
    .X(_03882_));
 sky130_fd_sc_hd__nand2_1 _10211_ (.A(net8),
    .B(net54),
    .Y(_03883_));
 sky130_fd_sc_hd__xnor2_1 _10212_ (.A(_03882_),
    .B(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__a31o_1 _10213_ (.A1(net7),
    .A2(net54),
    .A3(_03752_),
    .B1(_03751_),
    .X(_03885_));
 sky130_fd_sc_hd__nand2_1 _10214_ (.A(_03884_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__xor2_1 _10215_ (.A(_03884_),
    .B(_03885_),
    .X(_03888_));
 sky130_fd_sc_hd__and4b_1 _10216_ (.A_N(net6),
    .B(net7),
    .C(net56),
    .D(net57),
    .X(_03889_));
 sky130_fd_sc_hd__o2bb2a_1 _10217_ (.A1_N(net7),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net6),
    .X(_03890_));
 sky130_fd_sc_hd__nor2_1 _10218_ (.A(_03889_),
    .B(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__xnor2_1 _10219_ (.A(_03888_),
    .B(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__a21bo_1 _10220_ (.A1(_03759_),
    .A2(_03762_),
    .B1_N(_03758_),
    .X(_03893_));
 sky130_fd_sc_hd__and2b_1 _10221_ (.A_N(_03892_),
    .B(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__xor2_1 _10222_ (.A(_03892_),
    .B(_03893_),
    .X(_03895_));
 sky130_fd_sc_hd__inv_2 _10223_ (.A(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__and2_1 _10224_ (.A(_03760_),
    .B(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__xor2_1 _10225_ (.A(_03760_),
    .B(_03895_),
    .X(_03899_));
 sky130_fd_sc_hd__a21o_1 _10226_ (.A1(_03802_),
    .A2(_03810_),
    .B1(_03809_),
    .X(_03900_));
 sky130_fd_sc_hd__nand2_1 _10227_ (.A(_03774_),
    .B(_03777_),
    .Y(_03901_));
 sky130_fd_sc_hd__a31o_1 _10228_ (.A1(net14),
    .A2(net48),
    .A3(_03798_),
    .B1(_03797_),
    .X(_03902_));
 sky130_fd_sc_hd__nand4_1 _10229_ (.A(net13),
    .B(net14),
    .C(net49),
    .D(net50),
    .Y(_03903_));
 sky130_fd_sc_hd__a22o_1 _10230_ (.A1(net14),
    .A2(net49),
    .B1(net50),
    .B2(net13),
    .X(_03904_));
 sky130_fd_sc_hd__a22o_1 _10231_ (.A1(net11),
    .A2(net51),
    .B1(_03903_),
    .B2(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__nand4_1 _10232_ (.A(net11),
    .B(net51),
    .C(_03903_),
    .D(_03904_),
    .Y(_03906_));
 sky130_fd_sc_hd__nand3_1 _10233_ (.A(_03902_),
    .B(_03905_),
    .C(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__a21o_1 _10234_ (.A1(_03905_),
    .A2(_03906_),
    .B1(_03902_),
    .X(_03908_));
 sky130_fd_sc_hd__nand3_1 _10235_ (.A(_03901_),
    .B(_03907_),
    .C(_03908_),
    .Y(_03910_));
 sky130_fd_sc_hd__a21o_1 _10236_ (.A1(_03907_),
    .A2(_03908_),
    .B1(_03901_),
    .X(_03911_));
 sky130_fd_sc_hd__and3_1 _10237_ (.A(_03900_),
    .B(_03910_),
    .C(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__a21oi_1 _10238_ (.A1(_03910_),
    .A2(_03911_),
    .B1(_03900_),
    .Y(_03913_));
 sky130_fd_sc_hd__a211oi_2 _10239_ (.A1(_03779_),
    .A2(_03781_),
    .B1(_03912_),
    .C1(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__o211a_1 _10240_ (.A1(_03912_),
    .A2(_03913_),
    .B1(_03779_),
    .C1(_03781_),
    .X(_03915_));
 sky130_fd_sc_hd__a211oi_1 _10241_ (.A1(_03784_),
    .A2(_03786_),
    .B1(_03914_),
    .C1(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__o211a_1 _10242_ (.A1(_03914_),
    .A2(_03915_),
    .B1(_03784_),
    .C1(_03786_),
    .X(_03917_));
 sky130_fd_sc_hd__nor3_1 _10243_ (.A(_03899_),
    .B(_03916_),
    .C(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__o21a_1 _10244_ (.A1(_03916_),
    .A2(_03917_),
    .B1(_03899_),
    .X(_03919_));
 sky130_fd_sc_hd__a211oi_2 _10245_ (.A1(_03831_),
    .A2(_03834_),
    .B1(_03918_),
    .C1(_03919_),
    .Y(_03921_));
 sky130_fd_sc_hd__a211o_1 _10246_ (.A1(_03831_),
    .A2(_03834_),
    .B1(_03918_),
    .C1(_03919_),
    .X(_03922_));
 sky130_fd_sc_hd__o211ai_1 _10247_ (.A1(_03918_),
    .A2(_03919_),
    .B1(_03831_),
    .C1(_03834_),
    .Y(_03923_));
 sky130_fd_sc_hd__o211a_1 _10248_ (.A1(_03788_),
    .A2(_03791_),
    .B1(_03922_),
    .C1(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__a211oi_1 _10249_ (.A1(_03922_),
    .A2(_03923_),
    .B1(_03788_),
    .C1(_03791_),
    .Y(_03925_));
 sky130_fd_sc_hd__and4_1 _10250_ (.A(net46),
    .B(net47),
    .C(net16),
    .D(net17),
    .X(_03926_));
 sky130_fd_sc_hd__a22o_1 _10251_ (.A1(net47),
    .A2(net16),
    .B1(net17),
    .B2(net46),
    .X(_03927_));
 sky130_fd_sc_hd__and2b_1 _10252_ (.A_N(_03926_),
    .B(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__nand2_1 _10253_ (.A(net15),
    .B(net48),
    .Y(_03929_));
 sky130_fd_sc_hd__xnor2_1 _10254_ (.A(_03928_),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__nand4_1 _10255_ (.A(net42),
    .B(net43),
    .C(net19),
    .D(net20),
    .Y(_03932_));
 sky130_fd_sc_hd__a22o_1 _10256_ (.A1(net43),
    .A2(net19),
    .B1(net20),
    .B2(net42),
    .X(_03933_));
 sky130_fd_sc_hd__and2_1 _10257_ (.A(net45),
    .B(net18),
    .X(_03934_));
 sky130_fd_sc_hd__a21o_1 _10258_ (.A1(_03932_),
    .A2(_03933_),
    .B1(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__nand3_1 _10259_ (.A(_03932_),
    .B(_03933_),
    .C(_03934_),
    .Y(_03936_));
 sky130_fd_sc_hd__a21bo_1 _10260_ (.A1(_03804_),
    .A2(_03805_),
    .B1_N(_03803_),
    .X(_03937_));
 sky130_fd_sc_hd__and3_1 _10261_ (.A(_03935_),
    .B(_03936_),
    .C(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__a21o_1 _10262_ (.A1(_03935_),
    .A2(_03936_),
    .B1(_03937_),
    .X(_03939_));
 sky130_fd_sc_hd__and2b_1 _10263_ (.A_N(_03938_),
    .B(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__xnor2_1 _10264_ (.A(_03930_),
    .B(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__nand2_1 _10265_ (.A(_03816_),
    .B(_03819_),
    .Y(_03943_));
 sky130_fd_sc_hd__a31o_1 _10266_ (.A1(net38),
    .A2(net24),
    .A3(_03838_),
    .B1(_03837_),
    .X(_03944_));
 sky130_fd_sc_hd__nand4_1 _10267_ (.A(net39),
    .B(net40),
    .C(net22),
    .D(net24),
    .Y(_03945_));
 sky130_fd_sc_hd__a22o_1 _10268_ (.A1(net40),
    .A2(net22),
    .B1(net24),
    .B2(net39),
    .X(_03946_));
 sky130_fd_sc_hd__a22o_1 _10269_ (.A1(net41),
    .A2(net21),
    .B1(_03945_),
    .B2(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__nand4_1 _10270_ (.A(net41),
    .B(net21),
    .C(_03945_),
    .D(_03946_),
    .Y(_03948_));
 sky130_fd_sc_hd__nand3_1 _10271_ (.A(_03944_),
    .B(_03947_),
    .C(_03948_),
    .Y(_03949_));
 sky130_fd_sc_hd__a21o_1 _10272_ (.A1(_03947_),
    .A2(_03948_),
    .B1(_03944_),
    .X(_03950_));
 sky130_fd_sc_hd__nand3_1 _10273_ (.A(_03943_),
    .B(_03949_),
    .C(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__a21o_1 _10274_ (.A1(_03949_),
    .A2(_03950_),
    .B1(_03943_),
    .X(_03952_));
 sky130_fd_sc_hd__a21bo_1 _10275_ (.A1(_03814_),
    .A2(_03821_),
    .B1_N(_03820_),
    .X(_03954_));
 sky130_fd_sc_hd__and3_2 _10276_ (.A(_03951_),
    .B(_03952_),
    .C(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__a21oi_1 _10277_ (.A1(_03951_),
    .A2(_03952_),
    .B1(_03954_),
    .Y(_03956_));
 sky130_fd_sc_hd__or3_2 _10278_ (.A(_03941_),
    .B(_03955_),
    .C(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__inv_2 _10279_ (.A(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__o21ai_2 _10280_ (.A1(_03955_),
    .A2(_03956_),
    .B1(_03941_),
    .Y(_03959_));
 sky130_fd_sc_hd__o211ai_4 _10281_ (.A1(_03843_),
    .A2(_03846_),
    .B1(_03957_),
    .C1(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__a211o_1 _10282_ (.A1(_03957_),
    .A2(_03959_),
    .B1(_03843_),
    .C1(_03846_),
    .X(_03961_));
 sky130_fd_sc_hd__o211ai_2 _10283_ (.A1(_03826_),
    .A2(_03829_),
    .B1(_03960_),
    .C1(_03961_),
    .Y(_03962_));
 sky130_fd_sc_hd__a211o_1 _10284_ (.A1(_03960_),
    .A2(_03961_),
    .B1(_03826_),
    .C1(_03829_),
    .X(_03963_));
 sky130_fd_sc_hd__o21ai_1 _10285_ (.A1(_03718_),
    .A2(_03841_),
    .B1(_03591_),
    .Y(_03965_));
 sky130_fd_sc_hd__nand2_2 _10286_ (.A(net38),
    .B(net25),
    .Y(_03966_));
 sky130_fd_sc_hd__xor2_4 _10287_ (.A(_03839_),
    .B(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__xor2_2 _10288_ (.A(_03718_),
    .B(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__nand2_1 _10289_ (.A(_03442_),
    .B(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__xnor2_4 _10290_ (.A(_03441_),
    .B(_03968_),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_1 _10291_ (.A(_03965_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__xnor2_1 _10292_ (.A(_03965_),
    .B(_03970_),
    .Y(_03972_));
 sky130_fd_sc_hd__xnor2_1 _10293_ (.A(_03465_),
    .B(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__o21a_1 _10294_ (.A1(_03466_),
    .A2(_03847_),
    .B1(_03464_),
    .X(_03974_));
 sky130_fd_sc_hd__and2b_1 _10295_ (.A_N(_03974_),
    .B(_03973_),
    .X(_03976_));
 sky130_fd_sc_hd__xnor2_1 _10296_ (.A(_03973_),
    .B(_03974_),
    .Y(_03977_));
 sky130_fd_sc_hd__and3_1 _10297_ (.A(_03962_),
    .B(_03963_),
    .C(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__a21oi_1 _10298_ (.A1(_03962_),
    .A2(_03963_),
    .B1(_03977_),
    .Y(_03979_));
 sky130_fd_sc_hd__a211o_1 _10299_ (.A1(_03850_),
    .A2(_03852_),
    .B1(_03978_),
    .C1(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__o211ai_1 _10300_ (.A1(_03978_),
    .A2(_03979_),
    .B1(_03850_),
    .C1(_03852_),
    .Y(_03981_));
 sky130_fd_sc_hd__or4bb_2 _10301_ (.A(_03924_),
    .B(_03925_),
    .C_N(_03980_),
    .D_N(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__a2bb2o_1 _10302_ (.A1_N(_03924_),
    .A2_N(_03925_),
    .B1(_03980_),
    .B2(_03981_),
    .X(_03983_));
 sky130_fd_sc_hd__o211a_2 _10303_ (.A1(_03854_),
    .A2(_03858_),
    .B1(_03982_),
    .C1(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__a211oi_2 _10304_ (.A1(_03982_),
    .A2(_03983_),
    .B1(_03854_),
    .C1(_03858_),
    .Y(_03985_));
 sky130_fd_sc_hd__a211oi_4 _10305_ (.A1(_03793_),
    .A2(_03795_),
    .B1(_03984_),
    .C1(_03985_),
    .Y(_03987_));
 sky130_fd_sc_hd__o211a_1 _10306_ (.A1(_03984_),
    .A2(_03985_),
    .B1(_03793_),
    .C1(_03795_),
    .X(_03988_));
 sky130_fd_sc_hd__a211oi_2 _10307_ (.A1(_03860_),
    .A2(_03862_),
    .B1(_03987_),
    .C1(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__inv_2 _10308_ (.A(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__o211a_1 _10309_ (.A1(_03987_),
    .A2(_03988_),
    .B1(_03860_),
    .C1(_03862_),
    .X(_03991_));
 sky130_fd_sc_hd__a211o_1 _10310_ (.A1(_03765_),
    .A2(_03769_),
    .B1(_03989_),
    .C1(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__o211ai_1 _10311_ (.A1(_03989_),
    .A2(_03991_),
    .B1(_03765_),
    .C1(_03769_),
    .Y(_03993_));
 sky130_fd_sc_hd__nand2_2 _10312_ (.A(_03992_),
    .B(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__xnor2_2 _10313_ (.A(_03879_),
    .B(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__o21ai_1 _10314_ (.A1(_03868_),
    .A2(_03869_),
    .B1(_03876_),
    .Y(_03996_));
 sky130_fd_sc_hd__xnor2_1 _10315_ (.A(_03995_),
    .B(_03996_),
    .Y(net104));
 sky130_fd_sc_hd__or2_1 _10316_ (.A(_03916_),
    .B(_03918_),
    .X(_03998_));
 sky130_fd_sc_hd__and4_1 _10317_ (.A(net10),
    .B(net11),
    .C(net52),
    .D(net53),
    .X(_03999_));
 sky130_fd_sc_hd__a22o_1 _10318_ (.A1(net11),
    .A2(net52),
    .B1(net53),
    .B2(net10),
    .X(_04000_));
 sky130_fd_sc_hd__and2b_1 _10319_ (.A_N(_03999_),
    .B(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__nand2_1 _10320_ (.A(net9),
    .B(net54),
    .Y(_04002_));
 sky130_fd_sc_hd__xnor2_1 _10321_ (.A(_04001_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__a31o_1 _10322_ (.A1(net8),
    .A2(net54),
    .A3(_03881_),
    .B1(_03880_),
    .X(_04004_));
 sky130_fd_sc_hd__nand2_1 _10323_ (.A(_04003_),
    .B(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__xor2_1 _10324_ (.A(_04003_),
    .B(_04004_),
    .X(_04006_));
 sky130_fd_sc_hd__and4b_1 _10325_ (.A_N(net7),
    .B(net8),
    .C(net56),
    .D(net57),
    .X(_04008_));
 sky130_fd_sc_hd__o2bb2a_1 _10326_ (.A1_N(net8),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net7),
    .X(_04009_));
 sky130_fd_sc_hd__nor2_1 _10327_ (.A(_04008_),
    .B(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__xnor2_1 _10328_ (.A(_04006_),
    .B(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__a21bo_1 _10329_ (.A1(_03888_),
    .A2(_03891_),
    .B1_N(_03886_),
    .X(_04012_));
 sky130_fd_sc_hd__nand2b_1 _10330_ (.A_N(_04011_),
    .B(_04012_),
    .Y(_04013_));
 sky130_fd_sc_hd__xor2_1 _10331_ (.A(_04011_),
    .B(_04012_),
    .X(_04014_));
 sky130_fd_sc_hd__inv_2 _10332_ (.A(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__nand2_1 _10333_ (.A(_03889_),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__xor2_1 _10334_ (.A(_03889_),
    .B(_04014_),
    .X(_04017_));
 sky130_fd_sc_hd__a21o_1 _10335_ (.A1(_03930_),
    .A2(_03939_),
    .B1(_03938_),
    .X(_04019_));
 sky130_fd_sc_hd__nand2_1 _10336_ (.A(_03903_),
    .B(_03906_),
    .Y(_04020_));
 sky130_fd_sc_hd__a31o_1 _10337_ (.A1(net15),
    .A2(net48),
    .A3(_03927_),
    .B1(_03926_),
    .X(_04021_));
 sky130_fd_sc_hd__nand4_2 _10338_ (.A(net14),
    .B(net15),
    .C(net49),
    .D(net50),
    .Y(_04022_));
 sky130_fd_sc_hd__a22o_1 _10339_ (.A1(net15),
    .A2(net49),
    .B1(net50),
    .B2(net14),
    .X(_04023_));
 sky130_fd_sc_hd__a22o_1 _10340_ (.A1(net13),
    .A2(net51),
    .B1(_04022_),
    .B2(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__nand4_2 _10341_ (.A(net13),
    .B(net51),
    .C(_04022_),
    .D(_04023_),
    .Y(_04025_));
 sky130_fd_sc_hd__nand3_2 _10342_ (.A(_04021_),
    .B(_04024_),
    .C(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__a21o_1 _10343_ (.A1(_04024_),
    .A2(_04025_),
    .B1(_04021_),
    .X(_04027_));
 sky130_fd_sc_hd__nand3_2 _10344_ (.A(_04020_),
    .B(_04026_),
    .C(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__a21o_1 _10345_ (.A1(_04026_),
    .A2(_04027_),
    .B1(_04020_),
    .X(_04030_));
 sky130_fd_sc_hd__and3_1 _10346_ (.A(_04019_),
    .B(_04028_),
    .C(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__nand3_1 _10347_ (.A(_04019_),
    .B(_04028_),
    .C(_04030_),
    .Y(_04032_));
 sky130_fd_sc_hd__a21oi_1 _10348_ (.A1(_04028_),
    .A2(_04030_),
    .B1(_04019_),
    .Y(_04033_));
 sky130_fd_sc_hd__a211o_1 _10349_ (.A1(_03907_),
    .A2(_03910_),
    .B1(_04031_),
    .C1(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__o211ai_1 _10350_ (.A1(_04031_),
    .A2(_04033_),
    .B1(_03907_),
    .C1(_03910_),
    .Y(_04035_));
 sky130_fd_sc_hd__o211a_1 _10351_ (.A1(_03912_),
    .A2(_03914_),
    .B1(_04034_),
    .C1(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__a211oi_1 _10352_ (.A1(_04034_),
    .A2(_04035_),
    .B1(_03912_),
    .C1(_03914_),
    .Y(_04037_));
 sky130_fd_sc_hd__nor3_2 _10353_ (.A(_04017_),
    .B(_04036_),
    .C(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__o21a_1 _10354_ (.A1(_04036_),
    .A2(_04037_),
    .B1(_04017_),
    .X(_04039_));
 sky130_fd_sc_hd__a211o_1 _10355_ (.A1(_03960_),
    .A2(_03962_),
    .B1(_04038_),
    .C1(_04039_),
    .X(_04041_));
 sky130_fd_sc_hd__o211ai_2 _10356_ (.A1(_04038_),
    .A2(_04039_),
    .B1(_03960_),
    .C1(_03962_),
    .Y(_04042_));
 sky130_fd_sc_hd__nand3_2 _10357_ (.A(_03998_),
    .B(_04041_),
    .C(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__a21o_1 _10358_ (.A1(_04041_),
    .A2(_04042_),
    .B1(_03998_),
    .X(_04044_));
 sky130_fd_sc_hd__o21ai_4 _10359_ (.A1(_03718_),
    .A2(_03967_),
    .B1(_03591_),
    .Y(_04045_));
 sky130_fd_sc_hd__xor2_4 _10360_ (.A(_03970_),
    .B(_04045_),
    .X(_04046_));
 sky130_fd_sc_hd__or2_2 _10361_ (.A(_03465_),
    .B(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__xnor2_1 _10362_ (.A(_03466_),
    .B(_04046_),
    .Y(_04048_));
 sky130_fd_sc_hd__o21ai_1 _10363_ (.A1(_03466_),
    .A2(_03972_),
    .B1(_03464_),
    .Y(_04049_));
 sky130_fd_sc_hd__and2_1 _10364_ (.A(_04048_),
    .B(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__xor2_1 _10365_ (.A(_04048_),
    .B(_04049_),
    .X(_04052_));
 sky130_fd_sc_hd__and4_1 _10366_ (.A(net46),
    .B(net47),
    .C(net17),
    .D(net18),
    .X(_04053_));
 sky130_fd_sc_hd__a22o_1 _10367_ (.A1(net47),
    .A2(net17),
    .B1(net18),
    .B2(net46),
    .X(_04054_));
 sky130_fd_sc_hd__and2b_1 _10368_ (.A_N(_04053_),
    .B(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__nand2_1 _10369_ (.A(net16),
    .B(net48),
    .Y(_04056_));
 sky130_fd_sc_hd__xnor2_1 _10370_ (.A(_04055_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__nand4_1 _10371_ (.A(net42),
    .B(net43),
    .C(net20),
    .D(net21),
    .Y(_04058_));
 sky130_fd_sc_hd__a22o_1 _10372_ (.A1(net43),
    .A2(net20),
    .B1(net21),
    .B2(net42),
    .X(_04059_));
 sky130_fd_sc_hd__and2_1 _10373_ (.A(net45),
    .B(net19),
    .X(_04060_));
 sky130_fd_sc_hd__a21o_1 _10374_ (.A1(_04058_),
    .A2(_04059_),
    .B1(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__nand3_1 _10375_ (.A(_04058_),
    .B(_04059_),
    .C(_04060_),
    .Y(_04062_));
 sky130_fd_sc_hd__a21bo_1 _10376_ (.A1(_03933_),
    .A2(_03934_),
    .B1_N(_03932_),
    .X(_04063_));
 sky130_fd_sc_hd__and3_1 _10377_ (.A(_04061_),
    .B(_04062_),
    .C(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__a21o_1 _10378_ (.A1(_04061_),
    .A2(_04062_),
    .B1(_04063_),
    .X(_04065_));
 sky130_fd_sc_hd__and2b_1 _10379_ (.A_N(_04064_),
    .B(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__xor2_1 _10380_ (.A(_04057_),
    .B(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__nand2_1 _10381_ (.A(_03945_),
    .B(_03948_),
    .Y(_04068_));
 sky130_fd_sc_hd__a21o_1 _10382_ (.A1(net38),
    .A2(_03838_),
    .B1(_03837_),
    .X(_04069_));
 sky130_fd_sc_hd__nand4_1 _10383_ (.A(net39),
    .B(net40),
    .C(net24),
    .D(net25),
    .Y(_04070_));
 sky130_fd_sc_hd__a22o_1 _10384_ (.A1(net40),
    .A2(net24),
    .B1(net25),
    .B2(net39),
    .X(_04071_));
 sky130_fd_sc_hd__a22o_1 _10385_ (.A1(net41),
    .A2(net22),
    .B1(_04070_),
    .B2(_04071_),
    .X(_04073_));
 sky130_fd_sc_hd__nand4_1 _10386_ (.A(net41),
    .B(net22),
    .C(_04070_),
    .D(_04071_),
    .Y(_04074_));
 sky130_fd_sc_hd__nand3_1 _10387_ (.A(_04069_),
    .B(_04073_),
    .C(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__a21o_1 _10388_ (.A1(_04073_),
    .A2(_04074_),
    .B1(_04069_),
    .X(_04076_));
 sky130_fd_sc_hd__nand3_1 _10389_ (.A(_04068_),
    .B(_04075_),
    .C(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__a21o_1 _10390_ (.A1(_04075_),
    .A2(_04076_),
    .B1(_04068_),
    .X(_04078_));
 sky130_fd_sc_hd__a21bo_1 _10391_ (.A1(_03943_),
    .A2(_03950_),
    .B1_N(_03949_),
    .X(_04079_));
 sky130_fd_sc_hd__nand3_1 _10392_ (.A(_04077_),
    .B(_04078_),
    .C(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__a21o_1 _10393_ (.A1(_04077_),
    .A2(_04078_),
    .B1(_04079_),
    .X(_04081_));
 sky130_fd_sc_hd__and3_1 _10394_ (.A(_04067_),
    .B(_04080_),
    .C(_04081_),
    .X(_04082_));
 sky130_fd_sc_hd__a21oi_1 _10395_ (.A1(_04080_),
    .A2(_04081_),
    .B1(_04067_),
    .Y(_04084_));
 sky130_fd_sc_hd__a211o_2 _10396_ (.A1(_03969_),
    .A2(_03971_),
    .B1(_04082_),
    .C1(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__o211ai_2 _10397_ (.A1(_04082_),
    .A2(_04084_),
    .B1(_03969_),
    .C1(_03971_),
    .Y(_04086_));
 sky130_fd_sc_hd__o211ai_4 _10398_ (.A1(_03955_),
    .A2(_03958_),
    .B1(_04085_),
    .C1(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__a211o_1 _10399_ (.A1(_04085_),
    .A2(_04086_),
    .B1(_03955_),
    .C1(_03958_),
    .X(_04088_));
 sky130_fd_sc_hd__a21o_1 _10400_ (.A1(_04087_),
    .A2(_04088_),
    .B1(_04052_),
    .X(_04089_));
 sky130_fd_sc_hd__nand3_1 _10401_ (.A(_04052_),
    .B(_04087_),
    .C(_04088_),
    .Y(_04090_));
 sky130_fd_sc_hd__o211a_1 _10402_ (.A1(_03976_),
    .A2(_03978_),
    .B1(_04089_),
    .C1(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__o211ai_1 _10403_ (.A1(_03976_),
    .A2(_03978_),
    .B1(_04089_),
    .C1(_04090_),
    .Y(_04092_));
 sky130_fd_sc_hd__a211o_1 _10404_ (.A1(_04089_),
    .A2(_04090_),
    .B1(_03976_),
    .C1(_03978_),
    .X(_04093_));
 sky130_fd_sc_hd__and4_1 _10405_ (.A(_04043_),
    .B(_04044_),
    .C(_04092_),
    .D(_04093_),
    .X(_04095_));
 sky130_fd_sc_hd__a22oi_2 _10406_ (.A1(_04043_),
    .A2(_04044_),
    .B1(_04092_),
    .B2(_04093_),
    .Y(_04096_));
 sky130_fd_sc_hd__a211o_2 _10407_ (.A1(_03980_),
    .A2(_03982_),
    .B1(_04095_),
    .C1(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__o211ai_2 _10408_ (.A1(_04095_),
    .A2(_04096_),
    .B1(_03980_),
    .C1(_03982_),
    .Y(_04098_));
 sky130_fd_sc_hd__o211ai_4 _10409_ (.A1(_03921_),
    .A2(_03924_),
    .B1(_04097_),
    .C1(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__a211o_1 _10410_ (.A1(_04097_),
    .A2(_04098_),
    .B1(_03921_),
    .C1(_03924_),
    .X(_04100_));
 sky130_fd_sc_hd__o211ai_4 _10411_ (.A1(_03984_),
    .A2(_03987_),
    .B1(_04099_),
    .C1(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__a211o_1 _10412_ (.A1(_04099_),
    .A2(_04100_),
    .B1(_03984_),
    .C1(_03987_),
    .X(_04102_));
 sky130_fd_sc_hd__o211a_1 _10413_ (.A1(_03894_),
    .A2(_03897_),
    .B1(_04101_),
    .C1(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__o211ai_1 _10414_ (.A1(_03894_),
    .A2(_03897_),
    .B1(_04101_),
    .C1(_04102_),
    .Y(_04104_));
 sky130_fd_sc_hd__a211oi_1 _10415_ (.A1(_04101_),
    .A2(_04102_),
    .B1(_03894_),
    .C1(_03897_),
    .Y(_04106_));
 sky130_fd_sc_hd__a211oi_1 _10416_ (.A1(_03990_),
    .A2(_03992_),
    .B1(_04103_),
    .C1(_04106_),
    .Y(_04107_));
 sky130_fd_sc_hd__o211a_1 _10417_ (.A1(_04103_),
    .A2(_04106_),
    .B1(_03990_),
    .C1(_03992_),
    .X(_04108_));
 sky130_fd_sc_hd__or2_1 _10418_ (.A(_04107_),
    .B(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__a211o_1 _10419_ (.A1(_03879_),
    .A2(_03994_),
    .B1(_03868_),
    .C1(_03869_),
    .X(_04110_));
 sky130_fd_sc_hd__o21a_1 _10420_ (.A1(_03879_),
    .A2(_03994_),
    .B1(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__o31a_1 _10421_ (.A1(_03870_),
    .A2(_03875_),
    .A3(_03995_),
    .B1(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__xor2_1 _10422_ (.A(_04109_),
    .B(_04112_),
    .X(net105));
 sky130_fd_sc_hd__and2_2 _10423_ (.A(_03463_),
    .B(_04046_),
    .X(_04113_));
 sky130_fd_sc_hd__nand2_4 _10424_ (.A(_03463_),
    .B(_04046_),
    .Y(_04114_));
 sky130_fd_sc_hd__nor2_1 _10425_ (.A(_03463_),
    .B(_04047_),
    .Y(_04116_));
 sky130_fd_sc_hd__o21a_4 _10426_ (.A1(_03463_),
    .A2(_04047_),
    .B1(_04114_),
    .X(_04117_));
 sky130_fd_sc_hd__o21ai_4 _10427_ (.A1(_03463_),
    .A2(_04047_),
    .B1(_04114_),
    .Y(_04118_));
 sky130_fd_sc_hd__a31o_1 _10428_ (.A1(_04077_),
    .A2(_04078_),
    .A3(_04079_),
    .B1(_04082_),
    .X(_04119_));
 sky130_fd_sc_hd__a21bo_4 _10429_ (.A1(_03970_),
    .A2(_04045_),
    .B1_N(_03969_),
    .X(_04120_));
 sky130_fd_sc_hd__and4_1 _10430_ (.A(net46),
    .B(net47),
    .C(net18),
    .D(net19),
    .X(_04121_));
 sky130_fd_sc_hd__a22o_1 _10431_ (.A1(net47),
    .A2(net18),
    .B1(net19),
    .B2(net46),
    .X(_04122_));
 sky130_fd_sc_hd__and2b_1 _10432_ (.A_N(_04121_),
    .B(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__nand2_1 _10433_ (.A(net48),
    .B(net17),
    .Y(_04124_));
 sky130_fd_sc_hd__xnor2_1 _10434_ (.A(_04123_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand4_1 _10435_ (.A(net42),
    .B(net43),
    .C(net21),
    .D(net22),
    .Y(_04127_));
 sky130_fd_sc_hd__a22o_1 _10436_ (.A1(net43),
    .A2(net21),
    .B1(net22),
    .B2(net42),
    .X(_04128_));
 sky130_fd_sc_hd__and2_1 _10437_ (.A(net45),
    .B(net20),
    .X(_04129_));
 sky130_fd_sc_hd__a21o_1 _10438_ (.A1(_04127_),
    .A2(_04128_),
    .B1(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__nand3_1 _10439_ (.A(_04127_),
    .B(_04128_),
    .C(_04129_),
    .Y(_04131_));
 sky130_fd_sc_hd__a21bo_1 _10440_ (.A1(_04059_),
    .A2(_04060_),
    .B1_N(_04058_),
    .X(_04132_));
 sky130_fd_sc_hd__and3_1 _10441_ (.A(_04130_),
    .B(_04131_),
    .C(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__a21o_1 _10442_ (.A1(_04130_),
    .A2(_04131_),
    .B1(_04132_),
    .X(_04134_));
 sky130_fd_sc_hd__and2b_1 _10443_ (.A_N(_04133_),
    .B(_04134_),
    .X(_04135_));
 sky130_fd_sc_hd__xor2_1 _10444_ (.A(_04125_),
    .B(_04135_),
    .X(_04136_));
 sky130_fd_sc_hd__nand2_1 _10445_ (.A(_04070_),
    .B(_04074_),
    .Y(_04138_));
 sky130_fd_sc_hd__nand3_2 _10446_ (.A(net39),
    .B(net40),
    .C(net25),
    .Y(_04139_));
 sky130_fd_sc_hd__o21a_1 _10447_ (.A1(net39),
    .A2(net40),
    .B1(net25),
    .X(_04140_));
 sky130_fd_sc_hd__a22o_1 _10448_ (.A1(net41),
    .A2(net24),
    .B1(_04139_),
    .B2(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__nand4_1 _10449_ (.A(net41),
    .B(net24),
    .C(_04139_),
    .D(_04140_),
    .Y(_04142_));
 sky130_fd_sc_hd__nand3_1 _10450_ (.A(_04069_),
    .B(_04141_),
    .C(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__a21o_1 _10451_ (.A1(_04141_),
    .A2(_04142_),
    .B1(_04069_),
    .X(_04144_));
 sky130_fd_sc_hd__nand3_1 _10452_ (.A(_04138_),
    .B(_04143_),
    .C(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__a21o_1 _10453_ (.A1(_04143_),
    .A2(_04144_),
    .B1(_04138_),
    .X(_04146_));
 sky130_fd_sc_hd__a21bo_1 _10454_ (.A1(_04068_),
    .A2(_04076_),
    .B1_N(_04075_),
    .X(_04147_));
 sky130_fd_sc_hd__nand3_1 _10455_ (.A(_04145_),
    .B(_04146_),
    .C(_04147_),
    .Y(_04149_));
 sky130_fd_sc_hd__a21o_1 _10456_ (.A1(_04145_),
    .A2(_04146_),
    .B1(_04147_),
    .X(_04150_));
 sky130_fd_sc_hd__nand3_1 _10457_ (.A(_04136_),
    .B(_04149_),
    .C(_04150_),
    .Y(_04151_));
 sky130_fd_sc_hd__a21o_1 _10458_ (.A1(_04149_),
    .A2(_04150_),
    .B1(_04136_),
    .X(_04152_));
 sky130_fd_sc_hd__nand3_2 _10459_ (.A(_04120_),
    .B(_04151_),
    .C(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__a21o_1 _10460_ (.A1(_04151_),
    .A2(_04152_),
    .B1(_04120_),
    .X(_04154_));
 sky130_fd_sc_hd__nand3_2 _10461_ (.A(_04119_),
    .B(_04153_),
    .C(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__a21o_1 _10462_ (.A1(_04153_),
    .A2(_04154_),
    .B1(_04119_),
    .X(_04156_));
 sky130_fd_sc_hd__a21o_1 _10463_ (.A1(_04155_),
    .A2(_04156_),
    .B1(_04117_),
    .X(_04157_));
 sky130_fd_sc_hd__nand3_1 _10464_ (.A(_04117_),
    .B(_04155_),
    .C(_04156_),
    .Y(_04158_));
 sky130_fd_sc_hd__a31o_1 _10465_ (.A1(_04052_),
    .A2(_04087_),
    .A3(_04088_),
    .B1(_04050_),
    .X(_04160_));
 sky130_fd_sc_hd__and3_1 _10466_ (.A(_04157_),
    .B(_04158_),
    .C(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__nand3_1 _10467_ (.A(_04157_),
    .B(_04158_),
    .C(_04160_),
    .Y(_04162_));
 sky130_fd_sc_hd__a21oi_1 _10468_ (.A1(_04157_),
    .A2(_04158_),
    .B1(_04160_),
    .Y(_04163_));
 sky130_fd_sc_hd__and4_1 _10469_ (.A(net11),
    .B(net13),
    .C(net52),
    .D(net53),
    .X(_04164_));
 sky130_fd_sc_hd__a22o_1 _10470_ (.A1(net13),
    .A2(net52),
    .B1(net53),
    .B2(net11),
    .X(_04165_));
 sky130_fd_sc_hd__and2b_1 _10471_ (.A_N(_04164_),
    .B(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__nand2_1 _10472_ (.A(net10),
    .B(net54),
    .Y(_04167_));
 sky130_fd_sc_hd__xnor2_1 _10473_ (.A(_04166_),
    .B(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__a31o_1 _10474_ (.A1(net9),
    .A2(net54),
    .A3(_04000_),
    .B1(_03999_),
    .X(_04169_));
 sky130_fd_sc_hd__nand2_1 _10475_ (.A(_04168_),
    .B(_04169_),
    .Y(_04171_));
 sky130_fd_sc_hd__xor2_1 _10476_ (.A(_04168_),
    .B(_04169_),
    .X(_04172_));
 sky130_fd_sc_hd__and4b_1 _10477_ (.A_N(net8),
    .B(net9),
    .C(net56),
    .D(net57),
    .X(_04173_));
 sky130_fd_sc_hd__o2bb2a_1 _10478_ (.A1_N(net9),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net8),
    .X(_04174_));
 sky130_fd_sc_hd__nor2_1 _10479_ (.A(_04173_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__xnor2_1 _10480_ (.A(_04172_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__a21bo_1 _10481_ (.A1(_04006_),
    .A2(_04010_),
    .B1_N(_04005_),
    .X(_04177_));
 sky130_fd_sc_hd__and2b_1 _10482_ (.A_N(_04176_),
    .B(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__xor2_1 _10483_ (.A(_04176_),
    .B(_04177_),
    .X(_04179_));
 sky130_fd_sc_hd__inv_2 _10484_ (.A(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__xor2_1 _10485_ (.A(_04008_),
    .B(_04179_),
    .X(_04182_));
 sky130_fd_sc_hd__a21o_1 _10486_ (.A1(_04057_),
    .A2(_04065_),
    .B1(_04064_),
    .X(_04183_));
 sky130_fd_sc_hd__nand2_1 _10487_ (.A(_04022_),
    .B(_04025_),
    .Y(_04184_));
 sky130_fd_sc_hd__a31o_1 _10488_ (.A1(net16),
    .A2(net48),
    .A3(_04054_),
    .B1(_04053_),
    .X(_04185_));
 sky130_fd_sc_hd__nand4_1 _10489_ (.A(net15),
    .B(net16),
    .C(net49),
    .D(net50),
    .Y(_04186_));
 sky130_fd_sc_hd__a22o_1 _10490_ (.A1(net16),
    .A2(net49),
    .B1(net50),
    .B2(net15),
    .X(_04187_));
 sky130_fd_sc_hd__a22o_1 _10491_ (.A1(net14),
    .A2(net51),
    .B1(_04186_),
    .B2(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__nand4_1 _10492_ (.A(net14),
    .B(net51),
    .C(_04186_),
    .D(_04187_),
    .Y(_04189_));
 sky130_fd_sc_hd__nand3_1 _10493_ (.A(_04185_),
    .B(_04188_),
    .C(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__a21o_1 _10494_ (.A1(_04188_),
    .A2(_04189_),
    .B1(_04185_),
    .X(_04191_));
 sky130_fd_sc_hd__nand3_1 _10495_ (.A(_04184_),
    .B(_04190_),
    .C(_04191_),
    .Y(_04193_));
 sky130_fd_sc_hd__a21o_1 _10496_ (.A1(_04190_),
    .A2(_04191_),
    .B1(_04184_),
    .X(_04194_));
 sky130_fd_sc_hd__and3_1 _10497_ (.A(_04183_),
    .B(_04193_),
    .C(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__a21oi_1 _10498_ (.A1(_04193_),
    .A2(_04194_),
    .B1(_04183_),
    .Y(_04196_));
 sky130_fd_sc_hd__a211oi_2 _10499_ (.A1(_04026_),
    .A2(_04028_),
    .B1(_04195_),
    .C1(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__o211a_1 _10500_ (.A1(_04195_),
    .A2(_04196_),
    .B1(_04026_),
    .C1(_04028_),
    .X(_04198_));
 sky130_fd_sc_hd__a211oi_1 _10501_ (.A1(_04032_),
    .A2(_04034_),
    .B1(_04197_),
    .C1(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__o211a_1 _10502_ (.A1(_04197_),
    .A2(_04198_),
    .B1(_04032_),
    .C1(_04034_),
    .X(_04200_));
 sky130_fd_sc_hd__nor3_1 _10503_ (.A(_04182_),
    .B(_04199_),
    .C(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__o21a_1 _10504_ (.A1(_04199_),
    .A2(_04200_),
    .B1(_04182_),
    .X(_04202_));
 sky130_fd_sc_hd__a211o_1 _10505_ (.A1(_04085_),
    .A2(_04087_),
    .B1(_04201_),
    .C1(_04202_),
    .X(_04204_));
 sky130_fd_sc_hd__inv_2 _10506_ (.A(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__o211ai_1 _10507_ (.A1(_04201_),
    .A2(_04202_),
    .B1(_04085_),
    .C1(_04087_),
    .Y(_04206_));
 sky130_fd_sc_hd__o211a_1 _10508_ (.A1(_04036_),
    .A2(_04038_),
    .B1(_04204_),
    .C1(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__a211oi_1 _10509_ (.A1(_04204_),
    .A2(_04206_),
    .B1(_04036_),
    .C1(_04038_),
    .Y(_04208_));
 sky130_fd_sc_hd__or4_2 _10510_ (.A(_04161_),
    .B(_04163_),
    .C(_04207_),
    .D(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__o22ai_2 _10511_ (.A1(_04161_),
    .A2(_04163_),
    .B1(_04207_),
    .B2(_04208_),
    .Y(_04210_));
 sky130_fd_sc_hd__o211a_1 _10512_ (.A1(_04091_),
    .A2(_04095_),
    .B1(_04209_),
    .C1(_04210_),
    .X(_04211_));
 sky130_fd_sc_hd__a211oi_1 _10513_ (.A1(_04209_),
    .A2(_04210_),
    .B1(_04091_),
    .C1(_04095_),
    .Y(_04212_));
 sky130_fd_sc_hd__a211oi_2 _10514_ (.A1(_04041_),
    .A2(_04043_),
    .B1(_04211_),
    .C1(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__o211a_1 _10515_ (.A1(_04211_),
    .A2(_04212_),
    .B1(_04041_),
    .C1(_04043_),
    .X(_04215_));
 sky130_fd_sc_hd__a211oi_2 _10516_ (.A1(_04097_),
    .A2(_04099_),
    .B1(_04213_),
    .C1(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__o211a_1 _10517_ (.A1(_04213_),
    .A2(_04215_),
    .B1(_04097_),
    .C1(_04099_),
    .X(_04217_));
 sky130_fd_sc_hd__a211oi_2 _10518_ (.A1(_04013_),
    .A2(_04016_),
    .B1(_04216_),
    .C1(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__o211a_1 _10519_ (.A1(_04216_),
    .A2(_04217_),
    .B1(_04013_),
    .C1(_04016_),
    .X(_04219_));
 sky130_fd_sc_hd__o211a_1 _10520_ (.A1(_04218_),
    .A2(_04219_),
    .B1(_04101_),
    .C1(_04104_),
    .X(_04220_));
 sky130_fd_sc_hd__a211oi_1 _10521_ (.A1(_04101_),
    .A2(_04104_),
    .B1(_04218_),
    .C1(_04219_),
    .Y(_04221_));
 sky130_fd_sc_hd__nor2_1 _10522_ (.A(_04220_),
    .B(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__o21ba_1 _10523_ (.A1(_04109_),
    .A2(_04112_),
    .B1_N(_04107_),
    .X(_04223_));
 sky130_fd_sc_hd__xnor2_1 _10524_ (.A(_04222_),
    .B(_04223_),
    .Y(net106));
 sky130_fd_sc_hd__a21o_1 _10525_ (.A1(_04008_),
    .A2(_04180_),
    .B1(_04178_),
    .X(_04225_));
 sky130_fd_sc_hd__nand2_1 _10526_ (.A(_04149_),
    .B(_04151_),
    .Y(_04226_));
 sky130_fd_sc_hd__and4_1 _10527_ (.A(net46),
    .B(net47),
    .C(net19),
    .D(net20),
    .X(_04227_));
 sky130_fd_sc_hd__a22o_1 _10528_ (.A1(net47),
    .A2(net19),
    .B1(net20),
    .B2(net46),
    .X(_04228_));
 sky130_fd_sc_hd__and2b_1 _10529_ (.A_N(_04227_),
    .B(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__nand2_1 _10530_ (.A(net48),
    .B(net18),
    .Y(_04230_));
 sky130_fd_sc_hd__xnor2_1 _10531_ (.A(_04229_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand4_1 _10532_ (.A(net42),
    .B(net43),
    .C(net22),
    .D(net24),
    .Y(_04232_));
 sky130_fd_sc_hd__a22o_1 _10533_ (.A1(net43),
    .A2(net22),
    .B1(net24),
    .B2(net42),
    .X(_04233_));
 sky130_fd_sc_hd__and2_1 _10534_ (.A(net45),
    .B(net21),
    .X(_04234_));
 sky130_fd_sc_hd__a21o_1 _10535_ (.A1(_04232_),
    .A2(_04233_),
    .B1(_04234_),
    .X(_04236_));
 sky130_fd_sc_hd__nand3_1 _10536_ (.A(_04232_),
    .B(_04233_),
    .C(_04234_),
    .Y(_04237_));
 sky130_fd_sc_hd__a21bo_1 _10537_ (.A1(_04128_),
    .A2(_04129_),
    .B1_N(_04127_),
    .X(_04238_));
 sky130_fd_sc_hd__and3_1 _10538_ (.A(_04236_),
    .B(_04237_),
    .C(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__a21o_1 _10539_ (.A1(_04236_),
    .A2(_04237_),
    .B1(_04238_),
    .X(_04240_));
 sky130_fd_sc_hd__and2b_1 _10540_ (.A_N(_04239_),
    .B(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__xor2_1 _10541_ (.A(_04231_),
    .B(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__nand2_1 _10542_ (.A(_04139_),
    .B(_04142_),
    .Y(_04243_));
 sky130_fd_sc_hd__a22o_1 _10543_ (.A1(net41),
    .A2(net25),
    .B1(_04139_),
    .B2(_04140_),
    .X(_04244_));
 sky130_fd_sc_hd__nand3_1 _10544_ (.A(net41),
    .B(_04139_),
    .C(_04140_),
    .Y(_04245_));
 sky130_fd_sc_hd__nand3_2 _10545_ (.A(_04069_),
    .B(_04244_),
    .C(_04245_),
    .Y(_04247_));
 sky130_fd_sc_hd__a21o_1 _10546_ (.A1(_04244_),
    .A2(_04245_),
    .B1(_04069_),
    .X(_04248_));
 sky130_fd_sc_hd__nand3_1 _10547_ (.A(_04243_),
    .B(_04247_),
    .C(_04248_),
    .Y(_04249_));
 sky130_fd_sc_hd__a21o_1 _10548_ (.A1(_04247_),
    .A2(_04248_),
    .B1(_04243_),
    .X(_04250_));
 sky130_fd_sc_hd__a21bo_1 _10549_ (.A1(_04138_),
    .A2(_04144_),
    .B1_N(_04143_),
    .X(_04251_));
 sky130_fd_sc_hd__nand3_1 _10550_ (.A(_04249_),
    .B(_04250_),
    .C(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__a21o_1 _10551_ (.A1(_04249_),
    .A2(_04250_),
    .B1(_04251_),
    .X(_04253_));
 sky130_fd_sc_hd__nand3_1 _10552_ (.A(_04242_),
    .B(_04252_),
    .C(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__a21o_1 _10553_ (.A1(_04252_),
    .A2(_04253_),
    .B1(_04242_),
    .X(_04255_));
 sky130_fd_sc_hd__nand3_2 _10554_ (.A(_04120_),
    .B(_04254_),
    .C(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__a21o_1 _10555_ (.A1(_04254_),
    .A2(_04255_),
    .B1(_04120_),
    .X(_04258_));
 sky130_fd_sc_hd__nand3_2 _10556_ (.A(_04226_),
    .B(_04256_),
    .C(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__a21o_1 _10557_ (.A1(_04256_),
    .A2(_04258_),
    .B1(_04226_),
    .X(_04260_));
 sky130_fd_sc_hd__a21o_1 _10558_ (.A1(_04259_),
    .A2(_04260_),
    .B1(_04117_),
    .X(_04261_));
 sky130_fd_sc_hd__nand3_1 _10559_ (.A(_04117_),
    .B(_04259_),
    .C(_04260_),
    .Y(_04262_));
 sky130_fd_sc_hd__a31o_1 _10560_ (.A1(_04117_),
    .A2(_04155_),
    .A3(_04156_),
    .B1(_04113_),
    .X(_04263_));
 sky130_fd_sc_hd__and3_1 _10561_ (.A(_04261_),
    .B(_04262_),
    .C(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__inv_2 _10562_ (.A(_04264_),
    .Y(_04265_));
 sky130_fd_sc_hd__a21oi_1 _10563_ (.A1(_04261_),
    .A2(_04262_),
    .B1(_04263_),
    .Y(_04266_));
 sky130_fd_sc_hd__or2_1 _10564_ (.A(_04199_),
    .B(_04201_),
    .X(_04267_));
 sky130_fd_sc_hd__and4_1 _10565_ (.A(net13),
    .B(net14),
    .C(net52),
    .D(net53),
    .X(_04269_));
 sky130_fd_sc_hd__a22o_1 _10566_ (.A1(net14),
    .A2(net52),
    .B1(net53),
    .B2(net13),
    .X(_04270_));
 sky130_fd_sc_hd__and2b_1 _10567_ (.A_N(_04269_),
    .B(_04270_),
    .X(_04271_));
 sky130_fd_sc_hd__nand2_1 _10568_ (.A(net11),
    .B(net54),
    .Y(_04272_));
 sky130_fd_sc_hd__xnor2_1 _10569_ (.A(_04271_),
    .B(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__a31o_1 _10570_ (.A1(net10),
    .A2(net54),
    .A3(_04165_),
    .B1(_04164_),
    .X(_04274_));
 sky130_fd_sc_hd__nand2_1 _10571_ (.A(_04273_),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__xor2_1 _10572_ (.A(_04273_),
    .B(_04274_),
    .X(_04276_));
 sky130_fd_sc_hd__and4b_1 _10573_ (.A_N(net9),
    .B(net10),
    .C(net56),
    .D(net57),
    .X(_04277_));
 sky130_fd_sc_hd__o2bb2a_1 _10574_ (.A1_N(net10),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net9),
    .X(_04278_));
 sky130_fd_sc_hd__nor2_1 _10575_ (.A(_04277_),
    .B(_04278_),
    .Y(_04280_));
 sky130_fd_sc_hd__xnor2_1 _10576_ (.A(_04276_),
    .B(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__a21bo_1 _10577_ (.A1(_04172_),
    .A2(_04175_),
    .B1_N(_04171_),
    .X(_04282_));
 sky130_fd_sc_hd__nand2b_1 _10578_ (.A_N(_04281_),
    .B(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__xor2_1 _10579_ (.A(_04281_),
    .B(_04282_),
    .X(_04284_));
 sky130_fd_sc_hd__inv_2 _10580_ (.A(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__xor2_1 _10581_ (.A(_04173_),
    .B(_04284_),
    .X(_04286_));
 sky130_fd_sc_hd__a21o_1 _10582_ (.A1(_04125_),
    .A2(_04134_),
    .B1(_04133_),
    .X(_04287_));
 sky130_fd_sc_hd__nand2_1 _10583_ (.A(_04186_),
    .B(_04189_),
    .Y(_04288_));
 sky130_fd_sc_hd__a31o_1 _10584_ (.A1(net48),
    .A2(net17),
    .A3(_04122_),
    .B1(_04121_),
    .X(_04289_));
 sky130_fd_sc_hd__nand4_2 _10585_ (.A(net16),
    .B(net17),
    .C(net49),
    .D(net50),
    .Y(_04291_));
 sky130_fd_sc_hd__a22o_1 _10586_ (.A1(net17),
    .A2(net49),
    .B1(net50),
    .B2(net16),
    .X(_04292_));
 sky130_fd_sc_hd__a22o_1 _10587_ (.A1(net15),
    .A2(net51),
    .B1(_04291_),
    .B2(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__nand4_2 _10588_ (.A(net15),
    .B(net51),
    .C(_04291_),
    .D(_04292_),
    .Y(_04294_));
 sky130_fd_sc_hd__nand3_2 _10589_ (.A(_04289_),
    .B(_04293_),
    .C(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__a21o_1 _10590_ (.A1(_04293_),
    .A2(_04294_),
    .B1(_04289_),
    .X(_04296_));
 sky130_fd_sc_hd__nand3_2 _10591_ (.A(_04288_),
    .B(_04295_),
    .C(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__a21o_1 _10592_ (.A1(_04295_),
    .A2(_04296_),
    .B1(_04288_),
    .X(_04298_));
 sky130_fd_sc_hd__and3_1 _10593_ (.A(_04287_),
    .B(_04297_),
    .C(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__nand3_1 _10594_ (.A(_04287_),
    .B(_04297_),
    .C(_04298_),
    .Y(_04300_));
 sky130_fd_sc_hd__a21oi_1 _10595_ (.A1(_04297_),
    .A2(_04298_),
    .B1(_04287_),
    .Y(_04302_));
 sky130_fd_sc_hd__a211o_2 _10596_ (.A1(_04190_),
    .A2(_04193_),
    .B1(_04299_),
    .C1(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__o211ai_1 _10597_ (.A1(_04299_),
    .A2(_04302_),
    .B1(_04190_),
    .C1(_04193_),
    .Y(_04304_));
 sky130_fd_sc_hd__o211a_1 _10598_ (.A1(_04195_),
    .A2(_04197_),
    .B1(_04303_),
    .C1(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__a211oi_1 _10599_ (.A1(_04303_),
    .A2(_04304_),
    .B1(_04195_),
    .C1(_04197_),
    .Y(_04306_));
 sky130_fd_sc_hd__nor3_1 _10600_ (.A(_04286_),
    .B(_04305_),
    .C(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__o21a_1 _10601_ (.A1(_04305_),
    .A2(_04306_),
    .B1(_04286_),
    .X(_04308_));
 sky130_fd_sc_hd__a211o_1 _10602_ (.A1(_04153_),
    .A2(_04155_),
    .B1(_04307_),
    .C1(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__o211ai_1 _10603_ (.A1(_04307_),
    .A2(_04308_),
    .B1(_04153_),
    .C1(_04155_),
    .Y(_04310_));
 sky130_fd_sc_hd__and3_1 _10604_ (.A(_04267_),
    .B(_04309_),
    .C(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__inv_2 _10605_ (.A(_04311_),
    .Y(_04313_));
 sky130_fd_sc_hd__a21oi_1 _10606_ (.A1(_04309_),
    .A2(_04310_),
    .B1(_04267_),
    .Y(_04314_));
 sky130_fd_sc_hd__nor4_1 _10607_ (.A(_04264_),
    .B(_04266_),
    .C(_04311_),
    .D(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__or4_2 _10608_ (.A(_04264_),
    .B(_04266_),
    .C(_04311_),
    .D(_04314_),
    .X(_04316_));
 sky130_fd_sc_hd__o22a_1 _10609_ (.A1(_04264_),
    .A2(_04266_),
    .B1(_04311_),
    .B2(_04314_),
    .X(_04317_));
 sky130_fd_sc_hd__a211o_1 _10610_ (.A1(_04162_),
    .A2(_04209_),
    .B1(_04315_),
    .C1(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__o211ai_2 _10611_ (.A1(_04315_),
    .A2(_04317_),
    .B1(_04162_),
    .C1(_04209_),
    .Y(_04319_));
 sky130_fd_sc_hd__o211ai_2 _10612_ (.A1(_04205_),
    .A2(_04207_),
    .B1(_04318_),
    .C1(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__a211o_1 _10613_ (.A1(_04318_),
    .A2(_04319_),
    .B1(_04205_),
    .C1(_04207_),
    .X(_04321_));
 sky130_fd_sc_hd__o211a_1 _10614_ (.A1(_04211_),
    .A2(_04213_),
    .B1(_04320_),
    .C1(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__a211oi_1 _10615_ (.A1(_04320_),
    .A2(_04321_),
    .B1(_04211_),
    .C1(_04213_),
    .Y(_04324_));
 sky130_fd_sc_hd__nor2_1 _10616_ (.A(_04322_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__and2_1 _10617_ (.A(_04225_),
    .B(_04325_),
    .X(_04326_));
 sky130_fd_sc_hd__xnor2_1 _10618_ (.A(_04225_),
    .B(_04325_),
    .Y(_04327_));
 sky130_fd_sc_hd__or2_1 _10619_ (.A(_04216_),
    .B(_04218_),
    .X(_04328_));
 sky130_fd_sc_hd__and2b_1 _10620_ (.A_N(_04327_),
    .B(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__xnor2_1 _10621_ (.A(_04327_),
    .B(_04328_),
    .Y(_04330_));
 sky130_fd_sc_hd__or4_1 _10622_ (.A(_04107_),
    .B(_04108_),
    .C(_04220_),
    .D(_04221_),
    .X(_04331_));
 sky130_fd_sc_hd__nor3_1 _10623_ (.A(_03870_),
    .B(_03995_),
    .C(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__inv_2 _10624_ (.A(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__o21bai_1 _10625_ (.A1(_04107_),
    .A2(_04221_),
    .B1_N(_04220_),
    .Y(_04335_));
 sky130_fd_sc_hd__or2_1 _10626_ (.A(_04111_),
    .B(_04331_),
    .X(_04336_));
 sky130_fd_sc_hd__o211a_1 _10627_ (.A1(_03873_),
    .A2(_04333_),
    .B1(_04335_),
    .C1(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__o41a_2 _10628_ (.A1(_03344_),
    .A2(_03491_),
    .A3(_03871_),
    .A4(_04333_),
    .B1(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__and2_2 _10629_ (.A(_03348_),
    .B(_04337_),
    .X(_04339_));
 sky130_fd_sc_hd__a21oi_2 _10630_ (.A1(_03350_),
    .A2(_04339_),
    .B1(_04338_),
    .Y(_04340_));
 sky130_fd_sc_hd__xor2_1 _10631_ (.A(_04330_),
    .B(_04340_),
    .X(net107));
 sky130_fd_sc_hd__a21oi_1 _10632_ (.A1(_04330_),
    .A2(_04340_),
    .B1(_04329_),
    .Y(_04341_));
 sky130_fd_sc_hd__nand2_1 _10633_ (.A(_04252_),
    .B(_04254_),
    .Y(_04342_));
 sky130_fd_sc_hd__and4_1 _10634_ (.A(net46),
    .B(net47),
    .C(net20),
    .D(net21),
    .X(_04343_));
 sky130_fd_sc_hd__a22o_1 _10635_ (.A1(net47),
    .A2(net20),
    .B1(net21),
    .B2(net46),
    .X(_04345_));
 sky130_fd_sc_hd__and2b_1 _10636_ (.A_N(_04343_),
    .B(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _10637_ (.A(net48),
    .B(net19),
    .Y(_04347_));
 sky130_fd_sc_hd__xnor2_1 _10638_ (.A(_04346_),
    .B(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__and3_1 _10639_ (.A(net42),
    .B(net43),
    .C(net25),
    .X(_04349_));
 sky130_fd_sc_hd__nand4_1 _10640_ (.A(net42),
    .B(net43),
    .C(net24),
    .D(net25),
    .Y(_04350_));
 sky130_fd_sc_hd__a22o_1 _10641_ (.A1(net43),
    .A2(net24),
    .B1(net25),
    .B2(net42),
    .X(_04351_));
 sky130_fd_sc_hd__and2_1 _10642_ (.A(net45),
    .B(net22),
    .X(_04352_));
 sky130_fd_sc_hd__a21o_1 _10643_ (.A1(_04350_),
    .A2(_04351_),
    .B1(_04352_),
    .X(_04353_));
 sky130_fd_sc_hd__nand3_1 _10644_ (.A(_04350_),
    .B(_04351_),
    .C(_04352_),
    .Y(_04354_));
 sky130_fd_sc_hd__a21bo_1 _10645_ (.A1(_04233_),
    .A2(_04234_),
    .B1_N(_04232_),
    .X(_04356_));
 sky130_fd_sc_hd__and3_1 _10646_ (.A(_04353_),
    .B(_04354_),
    .C(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__a21o_1 _10647_ (.A1(_04353_),
    .A2(_04354_),
    .B1(_04356_),
    .X(_04358_));
 sky130_fd_sc_hd__nand2b_1 _10648_ (.A_N(_04357_),
    .B(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__xor2_1 _10649_ (.A(_04348_),
    .B(_04359_),
    .X(_04360_));
 sky130_fd_sc_hd__nand2_1 _10650_ (.A(_04139_),
    .B(_04245_),
    .Y(_04361_));
 sky130_fd_sc_hd__a21bo_1 _10651_ (.A1(_04247_),
    .A2(_04248_),
    .B1_N(_04361_),
    .X(_04362_));
 sky130_fd_sc_hd__nand3b_1 _10652_ (.A_N(_04361_),
    .B(_04248_),
    .C(_04247_),
    .Y(_04363_));
 sky130_fd_sc_hd__nor2_1 _10653_ (.A(_04139_),
    .B(_04247_),
    .Y(_04364_));
 sky130_fd_sc_hd__or2_2 _10654_ (.A(_04139_),
    .B(_04247_),
    .X(_04365_));
 sky130_fd_sc_hd__a41o_1 _10655_ (.A1(_04247_),
    .A2(_04249_),
    .A3(_04362_),
    .A4(_04363_),
    .B1(_04364_),
    .X(_04367_));
 sky130_fd_sc_hd__xor2_1 _10656_ (.A(_04360_),
    .B(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__nand2_1 _10657_ (.A(_04120_),
    .B(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__xnor2_1 _10658_ (.A(_04120_),
    .B(_04368_),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2b_1 _10659_ (.A_N(_04370_),
    .B(_04342_),
    .Y(_04371_));
 sky130_fd_sc_hd__xnor2_1 _10660_ (.A(_04342_),
    .B(_04370_),
    .Y(_04372_));
 sky130_fd_sc_hd__xnor2_1 _10661_ (.A(_04118_),
    .B(_04372_),
    .Y(_04373_));
 sky130_fd_sc_hd__a31o_1 _10662_ (.A1(_04117_),
    .A2(_04259_),
    .A3(_04260_),
    .B1(_04113_),
    .X(_04374_));
 sky130_fd_sc_hd__and2_1 _10663_ (.A(_04373_),
    .B(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__xor2_1 _10664_ (.A(_04373_),
    .B(_04374_),
    .X(_04376_));
 sky130_fd_sc_hd__and4_1 _10665_ (.A(net14),
    .B(net15),
    .C(net52),
    .D(net53),
    .X(_04378_));
 sky130_fd_sc_hd__a22o_1 _10666_ (.A1(net15),
    .A2(net52),
    .B1(net53),
    .B2(net14),
    .X(_04379_));
 sky130_fd_sc_hd__and2b_1 _10667_ (.A_N(_04378_),
    .B(_04379_),
    .X(_04380_));
 sky130_fd_sc_hd__nand2_1 _10668_ (.A(net13),
    .B(net54),
    .Y(_04381_));
 sky130_fd_sc_hd__xnor2_1 _10669_ (.A(_04380_),
    .B(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__a31o_1 _10670_ (.A1(net11),
    .A2(net54),
    .A3(_04270_),
    .B1(_04269_),
    .X(_04383_));
 sky130_fd_sc_hd__nand2_1 _10671_ (.A(_04382_),
    .B(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__xor2_1 _10672_ (.A(_04382_),
    .B(_04383_),
    .X(_04385_));
 sky130_fd_sc_hd__and4b_1 _10673_ (.A_N(net10),
    .B(net11),
    .C(net56),
    .D(net57),
    .X(_04386_));
 sky130_fd_sc_hd__o2bb2a_1 _10674_ (.A1_N(net11),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net10),
    .X(_04387_));
 sky130_fd_sc_hd__nor2_1 _10675_ (.A(_04386_),
    .B(_04387_),
    .Y(_04389_));
 sky130_fd_sc_hd__xnor2_1 _10676_ (.A(_04385_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__a21bo_1 _10677_ (.A1(_04276_),
    .A2(_04280_),
    .B1_N(_04275_),
    .X(_04391_));
 sky130_fd_sc_hd__and2b_1 _10678_ (.A_N(_04390_),
    .B(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__xor2_1 _10679_ (.A(_04390_),
    .B(_04391_),
    .X(_04393_));
 sky130_fd_sc_hd__inv_2 _10680_ (.A(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hd__and2_1 _10681_ (.A(_04277_),
    .B(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__xor2_1 _10682_ (.A(_04277_),
    .B(_04393_),
    .X(_04396_));
 sky130_fd_sc_hd__a21o_1 _10683_ (.A1(_04231_),
    .A2(_04240_),
    .B1(_04239_),
    .X(_04397_));
 sky130_fd_sc_hd__nand2_1 _10684_ (.A(_04291_),
    .B(_04294_),
    .Y(_04398_));
 sky130_fd_sc_hd__a31o_1 _10685_ (.A1(net48),
    .A2(net18),
    .A3(_04228_),
    .B1(_04227_),
    .X(_04400_));
 sky130_fd_sc_hd__nand4_2 _10686_ (.A(net17),
    .B(net49),
    .C(net18),
    .D(net50),
    .Y(_04401_));
 sky130_fd_sc_hd__a22o_1 _10687_ (.A1(net49),
    .A2(net18),
    .B1(net50),
    .B2(net17),
    .X(_04402_));
 sky130_fd_sc_hd__a22o_1 _10688_ (.A1(net16),
    .A2(net51),
    .B1(_04401_),
    .B2(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__nand4_2 _10689_ (.A(net16),
    .B(net51),
    .C(_04401_),
    .D(_04402_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand3_2 _10690_ (.A(_04400_),
    .B(_04403_),
    .C(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__a21o_1 _10691_ (.A1(_04403_),
    .A2(_04404_),
    .B1(_04400_),
    .X(_04406_));
 sky130_fd_sc_hd__nand3_2 _10692_ (.A(_04398_),
    .B(_04405_),
    .C(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__a21o_1 _10693_ (.A1(_04405_),
    .A2(_04406_),
    .B1(_04398_),
    .X(_04408_));
 sky130_fd_sc_hd__and3_2 _10694_ (.A(_04397_),
    .B(_04407_),
    .C(_04408_),
    .X(_04409_));
 sky130_fd_sc_hd__a21oi_2 _10695_ (.A1(_04407_),
    .A2(_04408_),
    .B1(_04397_),
    .Y(_04411_));
 sky130_fd_sc_hd__a211oi_4 _10696_ (.A1(_04295_),
    .A2(_04297_),
    .B1(_04409_),
    .C1(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__o211a_1 _10697_ (.A1(_04409_),
    .A2(_04411_),
    .B1(_04295_),
    .C1(_04297_),
    .X(_04413_));
 sky130_fd_sc_hd__a211oi_4 _10698_ (.A1(_04300_),
    .A2(_04303_),
    .B1(_04412_),
    .C1(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__o211a_1 _10699_ (.A1(_04412_),
    .A2(_04413_),
    .B1(_04300_),
    .C1(_04303_),
    .X(_04415_));
 sky130_fd_sc_hd__nor3_2 _10700_ (.A(_04396_),
    .B(_04414_),
    .C(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__o21a_1 _10701_ (.A1(_04414_),
    .A2(_04415_),
    .B1(_04396_),
    .X(_04417_));
 sky130_fd_sc_hd__a211o_1 _10702_ (.A1(_04256_),
    .A2(_04259_),
    .B1(_04416_),
    .C1(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__o211ai_2 _10703_ (.A1(_04416_),
    .A2(_04417_),
    .B1(_04256_),
    .C1(_04259_),
    .Y(_04419_));
 sky130_fd_sc_hd__o211ai_2 _10704_ (.A1(_04305_),
    .A2(_04307_),
    .B1(_04418_),
    .C1(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__a211o_1 _10705_ (.A1(_04418_),
    .A2(_04419_),
    .B1(_04305_),
    .C1(_04307_),
    .X(_04422_));
 sky130_fd_sc_hd__and3_2 _10706_ (.A(_04376_),
    .B(_04420_),
    .C(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__a21oi_2 _10707_ (.A1(_04420_),
    .A2(_04422_),
    .B1(_04376_),
    .Y(_04424_));
 sky130_fd_sc_hd__a211oi_4 _10708_ (.A1(_04265_),
    .A2(_04316_),
    .B1(_04423_),
    .C1(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__o211a_1 _10709_ (.A1(_04423_),
    .A2(_04424_),
    .B1(_04265_),
    .C1(_04316_),
    .X(_04426_));
 sky130_fd_sc_hd__a211oi_4 _10710_ (.A1(_04309_),
    .A2(_04313_),
    .B1(_04425_),
    .C1(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__o211a_1 _10711_ (.A1(_04425_),
    .A2(_04426_),
    .B1(_04309_),
    .C1(_04313_),
    .X(_04428_));
 sky130_fd_sc_hd__a211oi_1 _10712_ (.A1(_04318_),
    .A2(_04320_),
    .B1(_04427_),
    .C1(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__o211a_1 _10713_ (.A1(_04427_),
    .A2(_04428_),
    .B1(_04318_),
    .C1(_04320_),
    .X(_04430_));
 sky130_fd_sc_hd__inv_2 _10714_ (.A(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__or2_1 _10715_ (.A(_04429_),
    .B(_04430_),
    .X(_04433_));
 sky130_fd_sc_hd__a21bo_1 _10716_ (.A1(_04173_),
    .A2(_04285_),
    .B1_N(_04283_),
    .X(_04434_));
 sky130_fd_sc_hd__xnor2_1 _10717_ (.A(_04433_),
    .B(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__or3_1 _10718_ (.A(_04322_),
    .B(_04326_),
    .C(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__o21ai_1 _10719_ (.A1(_04322_),
    .A2(_04326_),
    .B1(_04435_),
    .Y(_04437_));
 sky130_fd_sc_hd__and2_1 _10720_ (.A(_04436_),
    .B(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__xnor2_1 _10721_ (.A(_04341_),
    .B(_04438_),
    .Y(net108));
 sky130_fd_sc_hd__o21a_1 _10722_ (.A1(_04360_),
    .A2(_04367_),
    .B1(_04365_),
    .X(_04439_));
 sky130_fd_sc_hd__and4_1 _10723_ (.A(net46),
    .B(net47),
    .C(net21),
    .D(net22),
    .X(_04440_));
 sky130_fd_sc_hd__a22o_1 _10724_ (.A1(net47),
    .A2(net21),
    .B1(net22),
    .B2(net46),
    .X(_04441_));
 sky130_fd_sc_hd__and2b_1 _10725_ (.A_N(_04440_),
    .B(_04441_),
    .X(_04443_));
 sky130_fd_sc_hd__nand2_1 _10726_ (.A(net48),
    .B(net20),
    .Y(_04444_));
 sky130_fd_sc_hd__xnor2_1 _10727_ (.A(_04443_),
    .B(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__o21ai_2 _10728_ (.A1(net42),
    .A2(net43),
    .B1(net25),
    .Y(_04446_));
 sky130_fd_sc_hd__nand2_1 _10729_ (.A(net45),
    .B(net24),
    .Y(_04447_));
 sky130_fd_sc_hd__o21ai_1 _10730_ (.A1(_04349_),
    .A2(_04446_),
    .B1(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__or3_1 _10731_ (.A(_04349_),
    .B(_04446_),
    .C(_04447_),
    .X(_04449_));
 sky130_fd_sc_hd__a21bo_1 _10732_ (.A1(_04351_),
    .A2(_04352_),
    .B1_N(_04350_),
    .X(_04450_));
 sky130_fd_sc_hd__and3_1 _10733_ (.A(_04448_),
    .B(_04449_),
    .C(_04450_),
    .X(_04451_));
 sky130_fd_sc_hd__a21o_1 _10734_ (.A1(_04448_),
    .A2(_04449_),
    .B1(_04450_),
    .X(_04452_));
 sky130_fd_sc_hd__and2b_1 _10735_ (.A_N(_04451_),
    .B(_04452_),
    .X(_04454_));
 sky130_fd_sc_hd__xnor2_1 _10736_ (.A(_04445_),
    .B(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__o21ai_4 _10737_ (.A1(_04248_),
    .A2(_04361_),
    .B1(_04365_),
    .Y(_04456_));
 sky130_fd_sc_hd__xor2_1 _10738_ (.A(_04455_),
    .B(_04456_),
    .X(_04457_));
 sky130_fd_sc_hd__and2_1 _10739_ (.A(_04120_),
    .B(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__xor2_1 _10740_ (.A(_04120_),
    .B(_04457_),
    .X(_04459_));
 sky130_fd_sc_hd__and2b_1 _10741_ (.A_N(_04439_),
    .B(_04459_),
    .X(_04460_));
 sky130_fd_sc_hd__xnor2_1 _10742_ (.A(_04439_),
    .B(_04459_),
    .Y(_04461_));
 sky130_fd_sc_hd__xnor2_1 _10743_ (.A(_04118_),
    .B(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__a21o_1 _10744_ (.A1(_04117_),
    .A2(_04372_),
    .B1(_04113_),
    .X(_04463_));
 sky130_fd_sc_hd__nand2_1 _10745_ (.A(_04462_),
    .B(_04463_),
    .Y(_04465_));
 sky130_fd_sc_hd__xor2_1 _10746_ (.A(_04462_),
    .B(_04463_),
    .X(_04466_));
 sky130_fd_sc_hd__and4_1 _10747_ (.A(net15),
    .B(net16),
    .C(net52),
    .D(net53),
    .X(_04467_));
 sky130_fd_sc_hd__a22o_1 _10748_ (.A1(net16),
    .A2(net52),
    .B1(net53),
    .B2(net15),
    .X(_04468_));
 sky130_fd_sc_hd__and2b_1 _10749_ (.A_N(_04467_),
    .B(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__nand2_1 _10750_ (.A(net14),
    .B(net54),
    .Y(_04470_));
 sky130_fd_sc_hd__xnor2_1 _10751_ (.A(_04469_),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__a31o_1 _10752_ (.A1(net13),
    .A2(net54),
    .A3(_04379_),
    .B1(_04378_),
    .X(_04472_));
 sky130_fd_sc_hd__nand2_1 _10753_ (.A(_04471_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__xor2_1 _10754_ (.A(_04471_),
    .B(_04472_),
    .X(_04474_));
 sky130_fd_sc_hd__and4b_1 _10755_ (.A_N(net11),
    .B(net13),
    .C(net56),
    .D(net57),
    .X(_04476_));
 sky130_fd_sc_hd__o2bb2a_1 _10756_ (.A1_N(net13),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net11),
    .X(_04477_));
 sky130_fd_sc_hd__nor2_1 _10757_ (.A(_04476_),
    .B(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__xnor2_1 _10758_ (.A(_04474_),
    .B(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__a21bo_1 _10759_ (.A1(_04385_),
    .A2(_04389_),
    .B1_N(_04384_),
    .X(_04480_));
 sky130_fd_sc_hd__nand2b_1 _10760_ (.A_N(_04479_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__xor2_1 _10761_ (.A(_04479_),
    .B(_04480_),
    .X(_04482_));
 sky130_fd_sc_hd__inv_2 _10762_ (.A(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__nand2_1 _10763_ (.A(_04386_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__xor2_1 _10764_ (.A(_04386_),
    .B(_04482_),
    .X(_04485_));
 sky130_fd_sc_hd__a21o_1 _10765_ (.A1(_04348_),
    .A2(_04358_),
    .B1(_04357_),
    .X(_04487_));
 sky130_fd_sc_hd__nand2_1 _10766_ (.A(_04401_),
    .B(_04404_),
    .Y(_04488_));
 sky130_fd_sc_hd__a31o_1 _10767_ (.A1(net48),
    .A2(net19),
    .A3(_04345_),
    .B1(_04343_),
    .X(_04489_));
 sky130_fd_sc_hd__nand4_2 _10768_ (.A(net49),
    .B(net18),
    .C(net50),
    .D(net19),
    .Y(_04490_));
 sky130_fd_sc_hd__a22o_1 _10769_ (.A1(net18),
    .A2(net50),
    .B1(net19),
    .B2(net49),
    .X(_04491_));
 sky130_fd_sc_hd__a22o_1 _10770_ (.A1(net17),
    .A2(net51),
    .B1(_04490_),
    .B2(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__nand4_2 _10771_ (.A(net17),
    .B(net51),
    .C(_04490_),
    .D(_04491_),
    .Y(_04493_));
 sky130_fd_sc_hd__nand3_2 _10772_ (.A(_04489_),
    .B(_04492_),
    .C(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__a21o_1 _10773_ (.A1(_04492_),
    .A2(_04493_),
    .B1(_04489_),
    .X(_04495_));
 sky130_fd_sc_hd__nand3_2 _10774_ (.A(_04488_),
    .B(_04494_),
    .C(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__a21o_1 _10775_ (.A1(_04494_),
    .A2(_04495_),
    .B1(_04488_),
    .X(_04498_));
 sky130_fd_sc_hd__and3_1 _10776_ (.A(_04487_),
    .B(_04496_),
    .C(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__nand3_1 _10777_ (.A(_04487_),
    .B(_04496_),
    .C(_04498_),
    .Y(_04500_));
 sky130_fd_sc_hd__a21oi_1 _10778_ (.A1(_04496_),
    .A2(_04498_),
    .B1(_04487_),
    .Y(_04501_));
 sky130_fd_sc_hd__a211o_2 _10779_ (.A1(_04405_),
    .A2(_04407_),
    .B1(_04499_),
    .C1(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__o211ai_1 _10780_ (.A1(_04499_),
    .A2(_04501_),
    .B1(_04405_),
    .C1(_04407_),
    .Y(_04503_));
 sky130_fd_sc_hd__o211a_1 _10781_ (.A1(_04409_),
    .A2(_04412_),
    .B1(_04502_),
    .C1(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__a211oi_1 _10782_ (.A1(_04502_),
    .A2(_04503_),
    .B1(_04409_),
    .C1(_04412_),
    .Y(_04505_));
 sky130_fd_sc_hd__nor3_2 _10783_ (.A(_04485_),
    .B(_04504_),
    .C(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__o21a_1 _10784_ (.A1(_04504_),
    .A2(_04505_),
    .B1(_04485_),
    .X(_04507_));
 sky130_fd_sc_hd__a211o_2 _10785_ (.A1(_04369_),
    .A2(_04371_),
    .B1(_04506_),
    .C1(_04507_),
    .X(_04509_));
 sky130_fd_sc_hd__o211ai_2 _10786_ (.A1(_04506_),
    .A2(_04507_),
    .B1(_04369_),
    .C1(_04371_),
    .Y(_04510_));
 sky130_fd_sc_hd__o211ai_4 _10787_ (.A1(_04414_),
    .A2(_04416_),
    .B1(_04509_),
    .C1(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__a211o_1 _10788_ (.A1(_04509_),
    .A2(_04510_),
    .B1(_04414_),
    .C1(_04416_),
    .X(_04512_));
 sky130_fd_sc_hd__nand3_2 _10789_ (.A(_04466_),
    .B(_04511_),
    .C(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__a21o_1 _10790_ (.A1(_04511_),
    .A2(_04512_),
    .B1(_04466_),
    .X(_04514_));
 sky130_fd_sc_hd__o211ai_2 _10791_ (.A1(_04375_),
    .A2(_04423_),
    .B1(_04513_),
    .C1(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__a211o_1 _10792_ (.A1(_04513_),
    .A2(_04514_),
    .B1(_04375_),
    .C1(_04423_),
    .X(_04516_));
 sky130_fd_sc_hd__nand2_1 _10793_ (.A(_04418_),
    .B(_04420_),
    .Y(_04517_));
 sky130_fd_sc_hd__nand3_2 _10794_ (.A(_04515_),
    .B(_04516_),
    .C(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__a21o_1 _10795_ (.A1(_04515_),
    .A2(_04516_),
    .B1(_04517_),
    .X(_04520_));
 sky130_fd_sc_hd__o211ai_4 _10796_ (.A1(_04425_),
    .A2(_04427_),
    .B1(_04518_),
    .C1(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__a211o_1 _10797_ (.A1(_04518_),
    .A2(_04520_),
    .B1(_04425_),
    .C1(_04427_),
    .X(_04522_));
 sky130_fd_sc_hd__o211ai_2 _10798_ (.A1(_04392_),
    .A2(_04395_),
    .B1(_04521_),
    .C1(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__a211o_1 _10799_ (.A1(_04521_),
    .A2(_04522_),
    .B1(_04392_),
    .C1(_04395_),
    .X(_04524_));
 sky130_fd_sc_hd__nand2_1 _10800_ (.A(_04523_),
    .B(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__a21oi_1 _10801_ (.A1(_04431_),
    .A2(_04434_),
    .B1(_04429_),
    .Y(_04526_));
 sky130_fd_sc_hd__nor2_1 _10802_ (.A(_04525_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__and2_1 _10803_ (.A(_04525_),
    .B(_04526_),
    .X(_04528_));
 sky130_fd_sc_hd__nor2_1 _10804_ (.A(_04527_),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__a21boi_1 _10805_ (.A1(_04329_),
    .A2(_04436_),
    .B1_N(_04437_),
    .Y(_04531_));
 sky130_fd_sc_hd__nand2_1 _10806_ (.A(_04330_),
    .B(_04438_),
    .Y(_04532_));
 sky130_fd_sc_hd__inv_2 _10807_ (.A(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__a21bo_1 _10808_ (.A1(_04340_),
    .A2(_04533_),
    .B1_N(_04531_),
    .X(_04534_));
 sky130_fd_sc_hd__xor2_1 _10809_ (.A(_04529_),
    .B(_04534_),
    .X(net110));
 sky130_fd_sc_hd__o21ai_1 _10810_ (.A1(_04455_),
    .A2(_04456_),
    .B1(_04365_),
    .Y(_04535_));
 sky130_fd_sc_hd__and4_1 _10811_ (.A(net46),
    .B(net47),
    .C(net22),
    .D(net24),
    .X(_04536_));
 sky130_fd_sc_hd__a22oi_1 _10812_ (.A1(net47),
    .A2(net22),
    .B1(net24),
    .B2(net46),
    .Y(_04537_));
 sky130_fd_sc_hd__nor2_1 _10813_ (.A(_04536_),
    .B(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__nand2_1 _10814_ (.A(net48),
    .B(net21),
    .Y(_04539_));
 sky130_fd_sc_hd__xnor2_1 _10815_ (.A(_04538_),
    .B(_04539_),
    .Y(_04541_));
 sky130_fd_sc_hd__o21bai_1 _10816_ (.A1(_04446_),
    .A2(_04447_),
    .B1_N(_04349_),
    .Y(_04542_));
 sky130_fd_sc_hd__nand2_1 _10817_ (.A(net45),
    .B(net25),
    .Y(_04543_));
 sky130_fd_sc_hd__o21ai_1 _10818_ (.A1(_04349_),
    .A2(_04446_),
    .B1(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__or3_1 _10819_ (.A(_04349_),
    .B(_04446_),
    .C(_04543_),
    .X(_04545_));
 sky130_fd_sc_hd__and2_1 _10820_ (.A(net45),
    .B(_04349_),
    .X(_04546_));
 sky130_fd_sc_hd__a21oi_1 _10821_ (.A1(_04544_),
    .A2(_04545_),
    .B1(_04542_),
    .Y(_04547_));
 sky130_fd_sc_hd__nor2_1 _10822_ (.A(_04546_),
    .B(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__xnor2_1 _10823_ (.A(_04541_),
    .B(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__xor2_1 _10824_ (.A(_04456_),
    .B(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__nand2_1 _10825_ (.A(_04120_),
    .B(_04550_),
    .Y(_04552_));
 sky130_fd_sc_hd__xnor2_1 _10826_ (.A(_04120_),
    .B(_04550_),
    .Y(_04553_));
 sky130_fd_sc_hd__nand2b_1 _10827_ (.A_N(_04553_),
    .B(_04535_),
    .Y(_04554_));
 sky130_fd_sc_hd__xor2_1 _10828_ (.A(_04535_),
    .B(_04553_),
    .X(_04555_));
 sky130_fd_sc_hd__and2_1 _10829_ (.A(_04118_),
    .B(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__nor2_1 _10830_ (.A(_04118_),
    .B(_04555_),
    .Y(_04557_));
 sky130_fd_sc_hd__or2_1 _10831_ (.A(_04556_),
    .B(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__a21oi_1 _10832_ (.A1(_04117_),
    .A2(_04461_),
    .B1(_04113_),
    .Y(_04559_));
 sky130_fd_sc_hd__nor2_1 _10833_ (.A(_04558_),
    .B(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__xor2_1 _10834_ (.A(_04558_),
    .B(_04559_),
    .X(_04561_));
 sky130_fd_sc_hd__and4_1 _10835_ (.A(net16),
    .B(net17),
    .C(net52),
    .D(net53),
    .X(_04563_));
 sky130_fd_sc_hd__a22oi_1 _10836_ (.A1(net17),
    .A2(net52),
    .B1(net53),
    .B2(net16),
    .Y(_04564_));
 sky130_fd_sc_hd__nor2_1 _10837_ (.A(_04563_),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_1 _10838_ (.A(net15),
    .B(net54),
    .Y(_04566_));
 sky130_fd_sc_hd__xnor2_1 _10839_ (.A(_04565_),
    .B(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__a31o_1 _10840_ (.A1(net14),
    .A2(net54),
    .A3(_04468_),
    .B1(_04467_),
    .X(_04568_));
 sky130_fd_sc_hd__nor2_1 _10841_ (.A(_04567_),
    .B(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__nand2_1 _10842_ (.A(_04567_),
    .B(_04568_),
    .Y(_04570_));
 sky130_fd_sc_hd__and2b_1 _10843_ (.A_N(_04569_),
    .B(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__and4b_1 _10844_ (.A_N(net13),
    .B(net14),
    .C(net56),
    .D(net57),
    .X(_04572_));
 sky130_fd_sc_hd__o2bb2a_1 _10845_ (.A1_N(net14),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net13),
    .X(_04574_));
 sky130_fd_sc_hd__nor2_1 _10846_ (.A(_04572_),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__xnor2_1 _10847_ (.A(_04571_),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__a21bo_1 _10848_ (.A1(_04474_),
    .A2(_04478_),
    .B1_N(_04473_),
    .X(_04577_));
 sky130_fd_sc_hd__and2b_1 _10849_ (.A_N(_04576_),
    .B(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__xor2_1 _10850_ (.A(_04576_),
    .B(_04577_),
    .X(_04579_));
 sky130_fd_sc_hd__inv_2 _10851_ (.A(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__xor2_1 _10852_ (.A(_04476_),
    .B(_04579_),
    .X(_04581_));
 sky130_fd_sc_hd__a21o_1 _10853_ (.A1(_04445_),
    .A2(_04452_),
    .B1(_04451_),
    .X(_04582_));
 sky130_fd_sc_hd__nand2_1 _10854_ (.A(_04490_),
    .B(_04493_),
    .Y(_04583_));
 sky130_fd_sc_hd__a31o_1 _10855_ (.A1(net48),
    .A2(net20),
    .A3(_04441_),
    .B1(_04440_),
    .X(_04585_));
 sky130_fd_sc_hd__nand4_1 _10856_ (.A(net49),
    .B(net50),
    .C(net19),
    .D(net20),
    .Y(_04586_));
 sky130_fd_sc_hd__a22o_1 _10857_ (.A1(net50),
    .A2(net19),
    .B1(net20),
    .B2(net49),
    .X(_04587_));
 sky130_fd_sc_hd__a22o_1 _10858_ (.A1(net18),
    .A2(net51),
    .B1(_04586_),
    .B2(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__nand4_1 _10859_ (.A(net18),
    .B(net51),
    .C(_04586_),
    .D(_04587_),
    .Y(_04589_));
 sky130_fd_sc_hd__nand3_1 _10860_ (.A(_04585_),
    .B(_04588_),
    .C(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__a21o_1 _10861_ (.A1(_04588_),
    .A2(_04589_),
    .B1(_04585_),
    .X(_04591_));
 sky130_fd_sc_hd__nand3_1 _10862_ (.A(_04583_),
    .B(_04590_),
    .C(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__a21o_1 _10863_ (.A1(_04590_),
    .A2(_04591_),
    .B1(_04583_),
    .X(_04593_));
 sky130_fd_sc_hd__and3_2 _10864_ (.A(_04582_),
    .B(_04592_),
    .C(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__a21oi_2 _10865_ (.A1(_04592_),
    .A2(_04593_),
    .B1(_04582_),
    .Y(_04596_));
 sky130_fd_sc_hd__a211oi_4 _10866_ (.A1(_04494_),
    .A2(_04496_),
    .B1(_04594_),
    .C1(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__o211a_1 _10867_ (.A1(_04594_),
    .A2(_04596_),
    .B1(_04494_),
    .C1(_04496_),
    .X(_04598_));
 sky130_fd_sc_hd__a211oi_4 _10868_ (.A1(_04500_),
    .A2(_04502_),
    .B1(_04597_),
    .C1(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__o211a_1 _10869_ (.A1(_04597_),
    .A2(_04598_),
    .B1(_04500_),
    .C1(_04502_),
    .X(_04600_));
 sky130_fd_sc_hd__or3_2 _10870_ (.A(_04581_),
    .B(_04599_),
    .C(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__inv_2 _10871_ (.A(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__o21ai_1 _10872_ (.A1(_04599_),
    .A2(_04600_),
    .B1(_04581_),
    .Y(_04603_));
 sky130_fd_sc_hd__o211ai_2 _10873_ (.A1(_04458_),
    .A2(_04460_),
    .B1(_04601_),
    .C1(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__a211o_1 _10874_ (.A1(_04601_),
    .A2(_04603_),
    .B1(_04458_),
    .C1(_04460_),
    .X(_04605_));
 sky130_fd_sc_hd__o211ai_2 _10875_ (.A1(_04504_),
    .A2(_04506_),
    .B1(_04604_),
    .C1(_04605_),
    .Y(_04607_));
 sky130_fd_sc_hd__a211o_1 _10876_ (.A1(_04604_),
    .A2(_04605_),
    .B1(_04504_),
    .C1(_04506_),
    .X(_04608_));
 sky130_fd_sc_hd__and3_1 _10877_ (.A(_04561_),
    .B(_04607_),
    .C(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__a21oi_1 _10878_ (.A1(_04607_),
    .A2(_04608_),
    .B1(_04561_),
    .Y(_04610_));
 sky130_fd_sc_hd__a211oi_2 _10879_ (.A1(_04465_),
    .A2(_04513_),
    .B1(_04609_),
    .C1(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__o211a_1 _10880_ (.A1(_04609_),
    .A2(_04610_),
    .B1(_04465_),
    .C1(_04513_),
    .X(_04612_));
 sky130_fd_sc_hd__a211oi_2 _10881_ (.A1(_04509_),
    .A2(_04511_),
    .B1(_04611_),
    .C1(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__o211a_1 _10882_ (.A1(_04611_),
    .A2(_04612_),
    .B1(_04509_),
    .C1(_04511_),
    .X(_04614_));
 sky130_fd_sc_hd__a211oi_1 _10883_ (.A1(_04515_),
    .A2(_04518_),
    .B1(_04613_),
    .C1(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__o211a_1 _10884_ (.A1(_04613_),
    .A2(_04614_),
    .B1(_04515_),
    .C1(_04518_),
    .X(_04616_));
 sky130_fd_sc_hd__a211oi_1 _10885_ (.A1(_04481_),
    .A2(_04484_),
    .B1(_04615_),
    .C1(_04616_),
    .Y(_04618_));
 sky130_fd_sc_hd__o211a_1 _10886_ (.A1(_04615_),
    .A2(_04616_),
    .B1(_04481_),
    .C1(_04484_),
    .X(_04619_));
 sky130_fd_sc_hd__o211a_1 _10887_ (.A1(_04618_),
    .A2(_04619_),
    .B1(_04521_),
    .C1(_04523_),
    .X(_04620_));
 sky130_fd_sc_hd__a211oi_1 _10888_ (.A1(_04521_),
    .A2(_04523_),
    .B1(_04618_),
    .C1(_04619_),
    .Y(_04621_));
 sky130_fd_sc_hd__nor2_1 _10889_ (.A(_04620_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__a21oi_1 _10890_ (.A1(_04529_),
    .A2(_04534_),
    .B1(_04527_),
    .Y(_04623_));
 sky130_fd_sc_hd__xnor2_1 _10891_ (.A(_04622_),
    .B(_04623_),
    .Y(net111));
 sky130_fd_sc_hd__o21ai_1 _10892_ (.A1(_04456_),
    .A2(_04549_),
    .B1(_04365_),
    .Y(_04624_));
 sky130_fd_sc_hd__and4_1 _10893_ (.A(net46),
    .B(net47),
    .C(net24),
    .D(net25),
    .X(_04625_));
 sky130_fd_sc_hd__a22oi_1 _10894_ (.A1(net47),
    .A2(net24),
    .B1(net25),
    .B2(net46),
    .Y(_04626_));
 sky130_fd_sc_hd__or2_1 _10895_ (.A(_04625_),
    .B(_04626_),
    .X(_04628_));
 sky130_fd_sc_hd__nand2_1 _10896_ (.A(net48),
    .B(net22),
    .Y(_04629_));
 sky130_fd_sc_hd__xnor2_1 _10897_ (.A(_04628_),
    .B(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__a21o_2 _10898_ (.A1(_04446_),
    .A2(_04543_),
    .B1(_04546_),
    .X(_04631_));
 sky130_fd_sc_hd__xnor2_1 _10899_ (.A(_04630_),
    .B(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__xor2_1 _10900_ (.A(_04456_),
    .B(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__and2_1 _10901_ (.A(_04120_),
    .B(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__xnor2_1 _10902_ (.A(_04120_),
    .B(_04633_),
    .Y(_04635_));
 sky130_fd_sc_hd__and2b_1 _10903_ (.A_N(_04635_),
    .B(_04624_),
    .X(_04636_));
 sky130_fd_sc_hd__xor2_1 _10904_ (.A(_04624_),
    .B(_04635_),
    .X(_04637_));
 sky130_fd_sc_hd__nor2_1 _10905_ (.A(_04118_),
    .B(_04637_),
    .Y(_04639_));
 sky130_fd_sc_hd__xnor2_1 _10906_ (.A(_04117_),
    .B(_04637_),
    .Y(_04640_));
 sky130_fd_sc_hd__o21ai_1 _10907_ (.A1(_04113_),
    .A2(_04557_),
    .B1(_04640_),
    .Y(_04641_));
 sky130_fd_sc_hd__or3_1 _10908_ (.A(_04113_),
    .B(_04557_),
    .C(_04640_),
    .X(_04642_));
 sky130_fd_sc_hd__and2_1 _10909_ (.A(_04641_),
    .B(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__and4_1 _10910_ (.A(net17),
    .B(net18),
    .C(net52),
    .D(net53),
    .X(_04644_));
 sky130_fd_sc_hd__a22oi_1 _10911_ (.A1(net18),
    .A2(net52),
    .B1(net53),
    .B2(net17),
    .Y(_04645_));
 sky130_fd_sc_hd__nor2_1 _10912_ (.A(_04644_),
    .B(_04645_),
    .Y(_04646_));
 sky130_fd_sc_hd__nand2_1 _10913_ (.A(net16),
    .B(net54),
    .Y(_04647_));
 sky130_fd_sc_hd__xnor2_1 _10914_ (.A(_04646_),
    .B(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__o21ba_1 _10915_ (.A1(_04564_),
    .A2(_04566_),
    .B1_N(_04563_),
    .X(_04650_));
 sky130_fd_sc_hd__nand2b_1 _10916_ (.A_N(_04650_),
    .B(_04648_),
    .Y(_04651_));
 sky130_fd_sc_hd__xnor2_1 _10917_ (.A(_04648_),
    .B(_04650_),
    .Y(_04652_));
 sky130_fd_sc_hd__and4b_1 _10918_ (.A_N(net14),
    .B(net15),
    .C(net56),
    .D(net57),
    .X(_04653_));
 sky130_fd_sc_hd__inv_2 _10919_ (.A(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__o2bb2a_1 _10920_ (.A1_N(net15),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net14),
    .X(_04655_));
 sky130_fd_sc_hd__nor2_1 _10921_ (.A(_04653_),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__or2_1 _10922_ (.A(_04652_),
    .B(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__nand2_1 _10923_ (.A(_04652_),
    .B(_04656_),
    .Y(_04658_));
 sky130_fd_sc_hd__nand2_1 _10924_ (.A(_04657_),
    .B(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__a21bo_1 _10925_ (.A1(_04571_),
    .A2(_04575_),
    .B1_N(_04570_),
    .X(_04661_));
 sky130_fd_sc_hd__nand2b_1 _10926_ (.A_N(_04659_),
    .B(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__xor2_1 _10927_ (.A(_04659_),
    .B(_04661_),
    .X(_04663_));
 sky130_fd_sc_hd__inv_2 _10928_ (.A(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__nand2_1 _10929_ (.A(_04572_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__xor2_1 _10930_ (.A(_04572_),
    .B(_04663_),
    .X(_04666_));
 sky130_fd_sc_hd__a21o_1 _10931_ (.A1(_04541_),
    .A2(_04548_),
    .B1(_04546_),
    .X(_04667_));
 sky130_fd_sc_hd__nand2_1 _10932_ (.A(_04586_),
    .B(_04589_),
    .Y(_04668_));
 sky130_fd_sc_hd__o21ba_1 _10933_ (.A1(_04537_),
    .A2(_04539_),
    .B1_N(_04536_),
    .X(_04669_));
 sky130_fd_sc_hd__and4_1 _10934_ (.A(net49),
    .B(net50),
    .C(net20),
    .D(net21),
    .X(_04670_));
 sky130_fd_sc_hd__a22oi_1 _10935_ (.A1(net50),
    .A2(net20),
    .B1(net21),
    .B2(net49),
    .Y(_04672_));
 sky130_fd_sc_hd__nor2_1 _10936_ (.A(_04670_),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__nand2_1 _10937_ (.A(net19),
    .B(net51),
    .Y(_04674_));
 sky130_fd_sc_hd__xnor2_1 _10938_ (.A(_04673_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__nand2b_1 _10939_ (.A_N(_04669_),
    .B(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__xnor2_1 _10940_ (.A(_04669_),
    .B(_04675_),
    .Y(_04677_));
 sky130_fd_sc_hd__nand2_1 _10941_ (.A(_04668_),
    .B(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hd__xor2_1 _10942_ (.A(_04668_),
    .B(_04677_),
    .X(_04679_));
 sky130_fd_sc_hd__nand2_1 _10943_ (.A(_04667_),
    .B(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__xnor2_1 _10944_ (.A(_04667_),
    .B(_04679_),
    .Y(_04681_));
 sky130_fd_sc_hd__a21o_1 _10945_ (.A1(_04590_),
    .A2(_04592_),
    .B1(_04681_),
    .X(_04683_));
 sky130_fd_sc_hd__nand3_1 _10946_ (.A(_04590_),
    .B(_04592_),
    .C(_04681_),
    .Y(_04684_));
 sky130_fd_sc_hd__o211a_1 _10947_ (.A1(_04594_),
    .A2(_04597_),
    .B1(_04683_),
    .C1(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__a211oi_1 _10948_ (.A1(_04683_),
    .A2(_04684_),
    .B1(_04594_),
    .C1(_04597_),
    .Y(_04686_));
 sky130_fd_sc_hd__nor3_2 _10949_ (.A(_04666_),
    .B(_04685_),
    .C(_04686_),
    .Y(_04687_));
 sky130_fd_sc_hd__o21a_1 _10950_ (.A1(_04685_),
    .A2(_04686_),
    .B1(_04666_),
    .X(_04688_));
 sky130_fd_sc_hd__a211o_2 _10951_ (.A1(_04552_),
    .A2(_04554_),
    .B1(_04687_),
    .C1(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__o211ai_2 _10952_ (.A1(_04687_),
    .A2(_04688_),
    .B1(_04552_),
    .C1(_04554_),
    .Y(_04690_));
 sky130_fd_sc_hd__o211ai_4 _10953_ (.A1(_04599_),
    .A2(_04602_),
    .B1(_04689_),
    .C1(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__a211o_1 _10954_ (.A1(_04689_),
    .A2(_04690_),
    .B1(_04599_),
    .C1(_04602_),
    .X(_04692_));
 sky130_fd_sc_hd__nand3_2 _10955_ (.A(_04643_),
    .B(_04691_),
    .C(_04692_),
    .Y(_04694_));
 sky130_fd_sc_hd__a21o_1 _10956_ (.A1(_04691_),
    .A2(_04692_),
    .B1(_04643_),
    .X(_04695_));
 sky130_fd_sc_hd__o211ai_2 _10957_ (.A1(_04560_),
    .A2(_04609_),
    .B1(_04694_),
    .C1(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__a211o_1 _10958_ (.A1(_04694_),
    .A2(_04695_),
    .B1(_04560_),
    .C1(_04609_),
    .X(_04697_));
 sky130_fd_sc_hd__nand2_1 _10959_ (.A(_04604_),
    .B(_04607_),
    .Y(_04698_));
 sky130_fd_sc_hd__nand3_1 _10960_ (.A(_04696_),
    .B(_04697_),
    .C(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hd__a21o_1 _10961_ (.A1(_04696_),
    .A2(_04697_),
    .B1(_04698_),
    .X(_04700_));
 sky130_fd_sc_hd__o211a_1 _10962_ (.A1(_04611_),
    .A2(_04613_),
    .B1(_04699_),
    .C1(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__a211o_1 _10963_ (.A1(_04699_),
    .A2(_04700_),
    .B1(_04611_),
    .C1(_04613_),
    .X(_04702_));
 sky130_fd_sc_hd__nand2b_1 _10964_ (.A_N(_04701_),
    .B(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__a21o_1 _10965_ (.A1(_04476_),
    .A2(_04580_),
    .B1(_04578_),
    .X(_04705_));
 sky130_fd_sc_hd__and3b_1 _10966_ (.A_N(_04701_),
    .B(_04702_),
    .C(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__xor2_1 _10967_ (.A(_04703_),
    .B(_04705_),
    .X(_04707_));
 sky130_fd_sc_hd__or2_1 _10968_ (.A(_04615_),
    .B(_04618_),
    .X(_04708_));
 sky130_fd_sc_hd__and2b_1 _10969_ (.A_N(_04707_),
    .B(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__xnor2_1 _10970_ (.A(_04707_),
    .B(_04708_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand2_1 _10971_ (.A(_04529_),
    .B(_04622_),
    .Y(_04711_));
 sky130_fd_sc_hd__nor2_1 _10972_ (.A(_04527_),
    .B(_04621_),
    .Y(_04712_));
 sky130_fd_sc_hd__o22ai_2 _10973_ (.A1(_04531_),
    .A2(_04711_),
    .B1(_04712_),
    .B2(_04620_),
    .Y(_04713_));
 sky130_fd_sc_hd__nor2_1 _10974_ (.A(_04532_),
    .B(_04711_),
    .Y(_04714_));
 sky130_fd_sc_hd__a21oi_1 _10975_ (.A1(_04340_),
    .A2(_04714_),
    .B1(_04713_),
    .Y(_04716_));
 sky130_fd_sc_hd__and2b_1 _10976_ (.A_N(_04716_),
    .B(_04710_),
    .X(_04717_));
 sky130_fd_sc_hd__and2b_1 _10977_ (.A_N(_04710_),
    .B(_04716_),
    .X(_04718_));
 sky130_fd_sc_hd__nor2_1 _10978_ (.A(_04717_),
    .B(_04718_),
    .Y(net112));
 sky130_fd_sc_hd__o21ai_1 _10979_ (.A1(_04456_),
    .A2(_04632_),
    .B1(_04365_),
    .Y(_04719_));
 sky130_fd_sc_hd__and3_1 _10980_ (.A(net46),
    .B(net47),
    .C(net25),
    .X(_04720_));
 sky130_fd_sc_hd__o21ai_1 _10981_ (.A1(net46),
    .A2(net47),
    .B1(net25),
    .Y(_04721_));
 sky130_fd_sc_hd__nor2_2 _10982_ (.A(_04720_),
    .B(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__nand2_1 _10983_ (.A(net48),
    .B(net24),
    .Y(_04723_));
 sky130_fd_sc_hd__xor2_1 _10984_ (.A(_04722_),
    .B(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__xor2_1 _10985_ (.A(_04631_),
    .B(_04724_),
    .X(_04726_));
 sky130_fd_sc_hd__nand2b_1 _10986_ (.A_N(_04456_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__xnor2_1 _10987_ (.A(_04456_),
    .B(_04726_),
    .Y(_04728_));
 sky130_fd_sc_hd__nand2_1 _10988_ (.A(_04120_),
    .B(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__xnor2_1 _10989_ (.A(_04120_),
    .B(_04728_),
    .Y(_04730_));
 sky130_fd_sc_hd__nand2b_1 _10990_ (.A_N(_04730_),
    .B(_04719_),
    .Y(_04731_));
 sky130_fd_sc_hd__xor2_1 _10991_ (.A(_04719_),
    .B(_04730_),
    .X(_04732_));
 sky130_fd_sc_hd__xnor2_1 _10992_ (.A(_04117_),
    .B(_04732_),
    .Y(_04733_));
 sky130_fd_sc_hd__o21a_1 _10993_ (.A1(_04113_),
    .A2(_04639_),
    .B1(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__nor3_1 _10994_ (.A(_04113_),
    .B(_04639_),
    .C(_04733_),
    .Y(_04735_));
 sky130_fd_sc_hd__nor2_1 _10995_ (.A(_04734_),
    .B(_04735_),
    .Y(_04737_));
 sky130_fd_sc_hd__and4_1 _10996_ (.A(net18),
    .B(net19),
    .C(net52),
    .D(net53),
    .X(_04738_));
 sky130_fd_sc_hd__a22oi_1 _10997_ (.A1(net19),
    .A2(net52),
    .B1(net53),
    .B2(net18),
    .Y(_04739_));
 sky130_fd_sc_hd__nor2_1 _10998_ (.A(_04738_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__nand2_1 _10999_ (.A(net17),
    .B(net54),
    .Y(_04741_));
 sky130_fd_sc_hd__xnor2_1 _11000_ (.A(_04740_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__o21ba_1 _11001_ (.A1(_04645_),
    .A2(_04647_),
    .B1_N(_04644_),
    .X(_04743_));
 sky130_fd_sc_hd__nand2b_1 _11002_ (.A_N(_04743_),
    .B(_04742_),
    .Y(_04744_));
 sky130_fd_sc_hd__xnor2_1 _11003_ (.A(_04742_),
    .B(_04743_),
    .Y(_04745_));
 sky130_fd_sc_hd__and4b_1 _11004_ (.A_N(net15),
    .B(net16),
    .C(net56),
    .D(net57),
    .X(_04746_));
 sky130_fd_sc_hd__o2bb2a_1 _11005_ (.A1_N(net16),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net15),
    .X(_04748_));
 sky130_fd_sc_hd__nor2_1 _11006_ (.A(_04746_),
    .B(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__or2_1 _11007_ (.A(_04745_),
    .B(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__nand2_1 _11008_ (.A(_04745_),
    .B(_04749_),
    .Y(_04751_));
 sky130_fd_sc_hd__nand2_1 _11009_ (.A(_04750_),
    .B(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__nand2_1 _11010_ (.A(_04651_),
    .B(_04658_),
    .Y(_04753_));
 sky130_fd_sc_hd__and2b_1 _11011_ (.A_N(_04752_),
    .B(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__xor2_1 _11012_ (.A(_04752_),
    .B(_04753_),
    .X(_04755_));
 sky130_fd_sc_hd__nor2_1 _11013_ (.A(_04654_),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__xnor2_1 _11014_ (.A(_04654_),
    .B(_04755_),
    .Y(_04757_));
 sky130_fd_sc_hd__o21bai_1 _11015_ (.A1(_04630_),
    .A2(_04631_),
    .B1_N(_04546_),
    .Y(_04759_));
 sky130_fd_sc_hd__o21ba_1 _11016_ (.A1(_04672_),
    .A2(_04674_),
    .B1_N(_04670_),
    .X(_04760_));
 sky130_fd_sc_hd__o21ba_1 _11017_ (.A1(_04626_),
    .A2(_04629_),
    .B1_N(_04625_),
    .X(_04761_));
 sky130_fd_sc_hd__and4_1 _11018_ (.A(net49),
    .B(net50),
    .C(net21),
    .D(net22),
    .X(_04762_));
 sky130_fd_sc_hd__a22oi_1 _11019_ (.A1(net50),
    .A2(net21),
    .B1(net22),
    .B2(net49),
    .Y(_04763_));
 sky130_fd_sc_hd__nor2_1 _11020_ (.A(_04762_),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__nand2_1 _11021_ (.A(net51),
    .B(net20),
    .Y(_04765_));
 sky130_fd_sc_hd__xnor2_1 _11022_ (.A(_04764_),
    .B(_04765_),
    .Y(_04766_));
 sky130_fd_sc_hd__nand2b_1 _11023_ (.A_N(_04761_),
    .B(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__xnor2_1 _11024_ (.A(_04761_),
    .B(_04766_),
    .Y(_04768_));
 sky130_fd_sc_hd__nand2b_1 _11025_ (.A_N(_04760_),
    .B(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__xnor2_1 _11026_ (.A(_04760_),
    .B(_04768_),
    .Y(_04770_));
 sky130_fd_sc_hd__and2_1 _11027_ (.A(_04759_),
    .B(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__xnor2_1 _11028_ (.A(_04759_),
    .B(_04770_),
    .Y(_04772_));
 sky130_fd_sc_hd__a21oi_2 _11029_ (.A1(_04676_),
    .A2(_04678_),
    .B1(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__and3_1 _11030_ (.A(_04676_),
    .B(_04678_),
    .C(_04772_),
    .X(_04774_));
 sky130_fd_sc_hd__a211oi_1 _11031_ (.A1(_04680_),
    .A2(_04683_),
    .B1(_04773_),
    .C1(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__a211o_1 _11032_ (.A1(_04680_),
    .A2(_04683_),
    .B1(_04773_),
    .C1(_04774_),
    .X(_04776_));
 sky130_fd_sc_hd__o211a_1 _11033_ (.A1(_04773_),
    .A2(_04774_),
    .B1(_04680_),
    .C1(_04683_),
    .X(_04777_));
 sky130_fd_sc_hd__or3_2 _11034_ (.A(_04757_),
    .B(_04775_),
    .C(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__o21ai_1 _11035_ (.A1(_04775_),
    .A2(_04777_),
    .B1(_04757_),
    .Y(_04780_));
 sky130_fd_sc_hd__o211ai_2 _11036_ (.A1(_04634_),
    .A2(_04636_),
    .B1(_04778_),
    .C1(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__a211o_1 _11037_ (.A1(_04778_),
    .A2(_04780_),
    .B1(_04634_),
    .C1(_04636_),
    .X(_04782_));
 sky130_fd_sc_hd__o211ai_2 _11038_ (.A1(_04685_),
    .A2(_04687_),
    .B1(_04781_),
    .C1(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__a211o_1 _11039_ (.A1(_04781_),
    .A2(_04782_),
    .B1(_04685_),
    .C1(_04687_),
    .X(_04784_));
 sky130_fd_sc_hd__and3_2 _11040_ (.A(_04737_),
    .B(_04783_),
    .C(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__a21oi_1 _11041_ (.A1(_04783_),
    .A2(_04784_),
    .B1(_04737_),
    .Y(_04786_));
 sky130_fd_sc_hd__a211oi_2 _11042_ (.A1(_04641_),
    .A2(_04694_),
    .B1(_04785_),
    .C1(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__o211a_1 _11043_ (.A1(_04785_),
    .A2(_04786_),
    .B1(_04641_),
    .C1(_04694_),
    .X(_04788_));
 sky130_fd_sc_hd__a211oi_2 _11044_ (.A1(_04689_),
    .A2(_04691_),
    .B1(_04787_),
    .C1(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__o211a_1 _11045_ (.A1(_04787_),
    .A2(_04788_),
    .B1(_04689_),
    .C1(_04691_),
    .X(_04791_));
 sky130_fd_sc_hd__a211oi_1 _11046_ (.A1(_04696_),
    .A2(_04699_),
    .B1(_04789_),
    .C1(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__o211a_1 _11047_ (.A1(_04789_),
    .A2(_04791_),
    .B1(_04696_),
    .C1(_04699_),
    .X(_04793_));
 sky130_fd_sc_hd__a211oi_1 _11048_ (.A1(_04662_),
    .A2(_04665_),
    .B1(_04792_),
    .C1(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__o211ai_1 _11049_ (.A1(_04792_),
    .A2(_04793_),
    .B1(_04662_),
    .C1(_04665_),
    .Y(_04795_));
 sky130_fd_sc_hd__and2b_1 _11050_ (.A_N(_04794_),
    .B(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__nor2_1 _11051_ (.A(_04701_),
    .B(_04706_),
    .Y(_04797_));
 sky130_fd_sc_hd__or3_1 _11052_ (.A(_04701_),
    .B(_04706_),
    .C(_04796_),
    .X(_04798_));
 sky130_fd_sc_hd__and2b_1 _11053_ (.A_N(_04797_),
    .B(_04796_),
    .X(_04799_));
 sky130_fd_sc_hd__xnor2_1 _11054_ (.A(_04796_),
    .B(_04797_),
    .Y(_04800_));
 sky130_fd_sc_hd__nor2_1 _11055_ (.A(_04709_),
    .B(_04717_),
    .Y(_04802_));
 sky130_fd_sc_hd__xnor2_1 _11056_ (.A(_04800_),
    .B(_04802_),
    .Y(net113));
 sky130_fd_sc_hd__nand2_1 _11057_ (.A(_04365_),
    .B(_04727_),
    .Y(_04803_));
 sky130_fd_sc_hd__a21o_1 _11058_ (.A1(net48),
    .A2(net25),
    .B1(_04722_),
    .X(_04804_));
 sky130_fd_sc_hd__a21bo_1 _11059_ (.A1(net48),
    .A2(_04722_),
    .B1_N(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__xor2_2 _11060_ (.A(_04631_),
    .B(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__and2b_1 _11061_ (.A_N(_04456_),
    .B(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__xnor2_2 _11062_ (.A(_04456_),
    .B(_04806_),
    .Y(_04808_));
 sky130_fd_sc_hd__and2_1 _11063_ (.A(_04120_),
    .B(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__xnor2_4 _11064_ (.A(_04120_),
    .B(_04808_),
    .Y(_04810_));
 sky130_fd_sc_hd__and2b_1 _11065_ (.A_N(_04810_),
    .B(_04803_),
    .X(_04812_));
 sky130_fd_sc_hd__xor2_1 _11066_ (.A(_04803_),
    .B(_04810_),
    .X(_04813_));
 sky130_fd_sc_hd__and2_1 _11067_ (.A(_04118_),
    .B(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__nor2_1 _11068_ (.A(_04118_),
    .B(_04813_),
    .Y(_04815_));
 sky130_fd_sc_hd__nor2_1 _11069_ (.A(_04814_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__o21a_1 _11070_ (.A1(_04118_),
    .A2(_04732_),
    .B1(_04114_),
    .X(_04817_));
 sky130_fd_sc_hd__or3_1 _11071_ (.A(_04814_),
    .B(_04815_),
    .C(_04817_),
    .X(_04818_));
 sky130_fd_sc_hd__xnor2_1 _11072_ (.A(_04816_),
    .B(_04817_),
    .Y(_04819_));
 sky130_fd_sc_hd__and4_1 _11073_ (.A(net19),
    .B(net20),
    .C(net52),
    .D(net53),
    .X(_04820_));
 sky130_fd_sc_hd__a22oi_1 _11074_ (.A1(net20),
    .A2(net52),
    .B1(net53),
    .B2(net19),
    .Y(_04821_));
 sky130_fd_sc_hd__nor2_1 _11075_ (.A(_04820_),
    .B(_04821_),
    .Y(_04823_));
 sky130_fd_sc_hd__nand2_1 _11076_ (.A(net18),
    .B(net54),
    .Y(_04824_));
 sky130_fd_sc_hd__xnor2_1 _11077_ (.A(_04823_),
    .B(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__o21ba_1 _11078_ (.A1(_04739_),
    .A2(_04741_),
    .B1_N(_04738_),
    .X(_04826_));
 sky130_fd_sc_hd__nand2b_1 _11079_ (.A_N(_04826_),
    .B(_04825_),
    .Y(_04827_));
 sky130_fd_sc_hd__xnor2_1 _11080_ (.A(_04825_),
    .B(_04826_),
    .Y(_04828_));
 sky130_fd_sc_hd__and4b_1 _11081_ (.A_N(net16),
    .B(net17),
    .C(net56),
    .D(net57),
    .X(_04829_));
 sky130_fd_sc_hd__inv_2 _11082_ (.A(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__o2bb2a_1 _11083_ (.A1_N(net17),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net16),
    .X(_04831_));
 sky130_fd_sc_hd__nor2_1 _11084_ (.A(_04829_),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__or2_1 _11085_ (.A(_04828_),
    .B(_04832_),
    .X(_04834_));
 sky130_fd_sc_hd__nand2_1 _11086_ (.A(_04828_),
    .B(_04832_),
    .Y(_04835_));
 sky130_fd_sc_hd__nand2_1 _11087_ (.A(_04834_),
    .B(_04835_),
    .Y(_04836_));
 sky130_fd_sc_hd__nand2_1 _11088_ (.A(_04744_),
    .B(_04751_),
    .Y(_04837_));
 sky130_fd_sc_hd__nand2b_1 _11089_ (.A_N(_04836_),
    .B(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__xor2_1 _11090_ (.A(_04836_),
    .B(_04837_),
    .X(_04839_));
 sky130_fd_sc_hd__inv_2 _11091_ (.A(_04839_),
    .Y(_04840_));
 sky130_fd_sc_hd__nand2_1 _11092_ (.A(_04746_),
    .B(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__xor2_1 _11093_ (.A(_04746_),
    .B(_04839_),
    .X(_04842_));
 sky130_fd_sc_hd__o21bai_1 _11094_ (.A1(_04631_),
    .A2(_04724_),
    .B1_N(_04546_),
    .Y(_04843_));
 sky130_fd_sc_hd__o21ba_1 _11095_ (.A1(_04763_),
    .A2(_04765_),
    .B1_N(_04762_),
    .X(_04845_));
 sky130_fd_sc_hd__o21ba_1 _11096_ (.A1(_04721_),
    .A2(_04723_),
    .B1_N(_04720_),
    .X(_04846_));
 sky130_fd_sc_hd__and4_1 _11097_ (.A(net49),
    .B(net50),
    .C(net22),
    .D(net24),
    .X(_04847_));
 sky130_fd_sc_hd__a22oi_1 _11098_ (.A1(net50),
    .A2(net22),
    .B1(net24),
    .B2(net49),
    .Y(_04848_));
 sky130_fd_sc_hd__nor2_1 _11099_ (.A(_04847_),
    .B(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__nand2_1 _11100_ (.A(net51),
    .B(net21),
    .Y(_04850_));
 sky130_fd_sc_hd__xnor2_1 _11101_ (.A(_04849_),
    .B(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__and2b_1 _11102_ (.A_N(_04846_),
    .B(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__xnor2_1 _11103_ (.A(_04846_),
    .B(_04851_),
    .Y(_04853_));
 sky130_fd_sc_hd__and2b_1 _11104_ (.A_N(_04845_),
    .B(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__xnor2_1 _11105_ (.A(_04845_),
    .B(_04853_),
    .Y(_04856_));
 sky130_fd_sc_hd__and2_1 _11106_ (.A(_04843_),
    .B(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__xnor2_1 _11107_ (.A(_04843_),
    .B(_04856_),
    .Y(_04858_));
 sky130_fd_sc_hd__a21oi_1 _11108_ (.A1(_04767_),
    .A2(_04769_),
    .B1(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__a21o_1 _11109_ (.A1(_04767_),
    .A2(_04769_),
    .B1(_04858_),
    .X(_04860_));
 sky130_fd_sc_hd__nand3_1 _11110_ (.A(_04767_),
    .B(_04769_),
    .C(_04858_),
    .Y(_04861_));
 sky130_fd_sc_hd__o211a_1 _11111_ (.A1(_04771_),
    .A2(_04773_),
    .B1(_04860_),
    .C1(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__a211oi_1 _11112_ (.A1(_04860_),
    .A2(_04861_),
    .B1(_04771_),
    .C1(_04773_),
    .Y(_04863_));
 sky130_fd_sc_hd__nor3_1 _11113_ (.A(_04842_),
    .B(_04862_),
    .C(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__o21a_1 _11114_ (.A1(_04862_),
    .A2(_04863_),
    .B1(_04842_),
    .X(_04865_));
 sky130_fd_sc_hd__a211oi_1 _11115_ (.A1(_04729_),
    .A2(_04731_),
    .B1(_04864_),
    .C1(_04865_),
    .Y(_04867_));
 sky130_fd_sc_hd__a211o_1 _11116_ (.A1(_04729_),
    .A2(_04731_),
    .B1(_04864_),
    .C1(_04865_),
    .X(_04868_));
 sky130_fd_sc_hd__o211a_1 _11117_ (.A1(_04864_),
    .A2(_04865_),
    .B1(_04729_),
    .C1(_04731_),
    .X(_04869_));
 sky130_fd_sc_hd__a211o_1 _11118_ (.A1(_04776_),
    .A2(_04778_),
    .B1(_04867_),
    .C1(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__o211ai_2 _11119_ (.A1(_04867_),
    .A2(_04869_),
    .B1(_04776_),
    .C1(_04778_),
    .Y(_04871_));
 sky130_fd_sc_hd__nand3_2 _11120_ (.A(_04819_),
    .B(_04870_),
    .C(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__a21o_1 _11121_ (.A1(_04870_),
    .A2(_04871_),
    .B1(_04819_),
    .X(_04873_));
 sky130_fd_sc_hd__o211ai_4 _11122_ (.A1(_04734_),
    .A2(_04785_),
    .B1(_04872_),
    .C1(_04873_),
    .Y(_04874_));
 sky130_fd_sc_hd__a211o_1 _11123_ (.A1(_04872_),
    .A2(_04873_),
    .B1(_04734_),
    .C1(_04785_),
    .X(_04875_));
 sky130_fd_sc_hd__nand2_1 _11124_ (.A(_04781_),
    .B(_04783_),
    .Y(_04876_));
 sky130_fd_sc_hd__nand3_2 _11125_ (.A(_04874_),
    .B(_04875_),
    .C(_04876_),
    .Y(_04878_));
 sky130_fd_sc_hd__a21o_1 _11126_ (.A1(_04874_),
    .A2(_04875_),
    .B1(_04876_),
    .X(_04879_));
 sky130_fd_sc_hd__o211ai_2 _11127_ (.A1(_04787_),
    .A2(_04789_),
    .B1(_04878_),
    .C1(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__a211o_1 _11128_ (.A1(_04878_),
    .A2(_04879_),
    .B1(_04787_),
    .C1(_04789_),
    .X(_04881_));
 sky130_fd_sc_hd__nand2_1 _11129_ (.A(_04880_),
    .B(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__nor2_1 _11130_ (.A(_04754_),
    .B(_04756_),
    .Y(_04883_));
 sky130_fd_sc_hd__o211ai_1 _11131_ (.A1(_04754_),
    .A2(_04756_),
    .B1(_04880_),
    .C1(_04881_),
    .Y(_04884_));
 sky130_fd_sc_hd__xnor2_1 _11132_ (.A(_04882_),
    .B(_04883_),
    .Y(_04885_));
 sky130_fd_sc_hd__or2_1 _11133_ (.A(_04792_),
    .B(_04794_),
    .X(_04886_));
 sky130_fd_sc_hd__and2b_1 _11134_ (.A_N(_04885_),
    .B(_04886_),
    .X(_04887_));
 sky130_fd_sc_hd__xnor2_1 _11135_ (.A(_04885_),
    .B(_04886_),
    .Y(_04889_));
 sky130_fd_sc_hd__a21oi_1 _11136_ (.A1(_04709_),
    .A2(_04798_),
    .B1(_04799_),
    .Y(_04890_));
 sky130_fd_sc_hd__nand2_1 _11137_ (.A(_04710_),
    .B(_04800_),
    .Y(_04891_));
 sky130_fd_sc_hd__o21ai_1 _11138_ (.A1(_04716_),
    .A2(_04891_),
    .B1(_04890_),
    .Y(_04892_));
 sky130_fd_sc_hd__xor2_1 _11139_ (.A(_04889_),
    .B(_04892_),
    .X(net114));
 sky130_fd_sc_hd__nor2_2 _11140_ (.A(_04364_),
    .B(_04807_),
    .Y(_04893_));
 sky130_fd_sc_hd__xnor2_4 _11141_ (.A(_04810_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__xnor2_1 _11142_ (.A(_04117_),
    .B(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__o21a_1 _11143_ (.A1(_04113_),
    .A2(_04815_),
    .B1(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__nor3_1 _11144_ (.A(_04113_),
    .B(_04815_),
    .C(_04895_),
    .Y(_04897_));
 sky130_fd_sc_hd__nor2_1 _11145_ (.A(_04896_),
    .B(_04897_),
    .Y(_04899_));
 sky130_fd_sc_hd__nor2_1 _11146_ (.A(_04862_),
    .B(_04864_),
    .Y(_04900_));
 sky130_fd_sc_hd__and4_1 _11147_ (.A(net20),
    .B(net52),
    .C(net21),
    .D(net53),
    .X(_04901_));
 sky130_fd_sc_hd__a22oi_1 _11148_ (.A1(net52),
    .A2(net21),
    .B1(net53),
    .B2(net20),
    .Y(_04902_));
 sky130_fd_sc_hd__nor2_1 _11149_ (.A(_04901_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__nand2_1 _11150_ (.A(net19),
    .B(net54),
    .Y(_04904_));
 sky130_fd_sc_hd__xnor2_1 _11151_ (.A(_04903_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__o21ba_1 _11152_ (.A1(_04821_),
    .A2(_04824_),
    .B1_N(_04820_),
    .X(_04906_));
 sky130_fd_sc_hd__nand2b_1 _11153_ (.A_N(_04906_),
    .B(_04905_),
    .Y(_04907_));
 sky130_fd_sc_hd__xnor2_1 _11154_ (.A(_04905_),
    .B(_04906_),
    .Y(_04908_));
 sky130_fd_sc_hd__and4b_1 _11155_ (.A_N(net17),
    .B(net18),
    .C(net56),
    .D(net57),
    .X(_04910_));
 sky130_fd_sc_hd__inv_2 _11156_ (.A(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__o2bb2a_1 _11157_ (.A1_N(net18),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net17),
    .X(_04912_));
 sky130_fd_sc_hd__nor2_1 _11158_ (.A(_04910_),
    .B(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__or2_1 _11159_ (.A(_04908_),
    .B(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__nand2_1 _11160_ (.A(_04908_),
    .B(_04913_),
    .Y(_04915_));
 sky130_fd_sc_hd__nand2_1 _11161_ (.A(_04914_),
    .B(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__nand2_1 _11162_ (.A(_04827_),
    .B(_04835_),
    .Y(_04917_));
 sky130_fd_sc_hd__and3_1 _11163_ (.A(_04914_),
    .B(_04915_),
    .C(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__xor2_1 _11164_ (.A(_04916_),
    .B(_04917_),
    .X(_04919_));
 sky130_fd_sc_hd__xnor2_1 _11165_ (.A(_04830_),
    .B(_04919_),
    .Y(_04921_));
 sky130_fd_sc_hd__nor2_1 _11166_ (.A(_04852_),
    .B(_04854_),
    .Y(_04922_));
 sky130_fd_sc_hd__o21ba_4 _11167_ (.A1(_04631_),
    .A2(_04805_),
    .B1_N(_04546_),
    .X(_04923_));
 sky130_fd_sc_hd__a31o_1 _11168_ (.A1(net51),
    .A2(net21),
    .A3(_04849_),
    .B1(_04847_),
    .X(_04924_));
 sky130_fd_sc_hd__a21oi_4 _11169_ (.A1(net48),
    .A2(_04722_),
    .B1(_04720_),
    .Y(_04925_));
 sky130_fd_sc_hd__and4_1 _11170_ (.A(net49),
    .B(net50),
    .C(net24),
    .D(net25),
    .X(_04926_));
 sky130_fd_sc_hd__a22oi_1 _11171_ (.A1(net50),
    .A2(net24),
    .B1(net25),
    .B2(net49),
    .Y(_04927_));
 sky130_fd_sc_hd__or2_1 _11172_ (.A(_04926_),
    .B(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__nand2_1 _11173_ (.A(net51),
    .B(net22),
    .Y(_04929_));
 sky130_fd_sc_hd__nor2_1 _11174_ (.A(_04928_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__xor2_1 _11175_ (.A(_04928_),
    .B(_04929_),
    .X(_04932_));
 sky130_fd_sc_hd__and2b_1 _11176_ (.A_N(_04925_),
    .B(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__xnor2_1 _11177_ (.A(_04925_),
    .B(_04932_),
    .Y(_04934_));
 sky130_fd_sc_hd__xnor2_1 _11178_ (.A(_04924_),
    .B(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__or2_1 _11179_ (.A(_04923_),
    .B(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__xor2_1 _11180_ (.A(_04923_),
    .B(_04935_),
    .X(_04937_));
 sky130_fd_sc_hd__nand2b_1 _11181_ (.A_N(_04922_),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__xnor2_1 _11182_ (.A(_04922_),
    .B(_04937_),
    .Y(_04939_));
 sky130_fd_sc_hd__o21a_1 _11183_ (.A1(_04857_),
    .A2(_04859_),
    .B1(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__nor3_1 _11184_ (.A(_04857_),
    .B(_04859_),
    .C(_04939_),
    .Y(_04941_));
 sky130_fd_sc_hd__or3_1 _11185_ (.A(_04921_),
    .B(_04940_),
    .C(_04941_),
    .X(_04943_));
 sky130_fd_sc_hd__o21ai_1 _11186_ (.A1(_04940_),
    .A2(_04941_),
    .B1(_04921_),
    .Y(_04944_));
 sky130_fd_sc_hd__o211ai_2 _11187_ (.A1(_04809_),
    .A2(_04812_),
    .B1(_04943_),
    .C1(_04944_),
    .Y(_04945_));
 sky130_fd_sc_hd__a211o_1 _11188_ (.A1(_04943_),
    .A2(_04944_),
    .B1(_04809_),
    .C1(_04812_),
    .X(_04946_));
 sky130_fd_sc_hd__nand3b_1 _11189_ (.A_N(_04900_),
    .B(_04945_),
    .C(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hd__a21bo_1 _11190_ (.A1(_04945_),
    .A2(_04946_),
    .B1_N(_04900_),
    .X(_04948_));
 sky130_fd_sc_hd__a21oi_1 _11191_ (.A1(_04947_),
    .A2(_04948_),
    .B1(_04899_),
    .Y(_04949_));
 sky130_fd_sc_hd__and3_1 _11192_ (.A(_04899_),
    .B(_04947_),
    .C(_04948_),
    .X(_04950_));
 sky130_fd_sc_hd__a211oi_2 _11193_ (.A1(_04818_),
    .A2(_04872_),
    .B1(_04949_),
    .C1(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__o211a_1 _11194_ (.A1(_04949_),
    .A2(_04950_),
    .B1(_04818_),
    .C1(_04872_),
    .X(_04952_));
 sky130_fd_sc_hd__a211oi_2 _11195_ (.A1(_04868_),
    .A2(_04870_),
    .B1(_04951_),
    .C1(_04952_),
    .Y(_04954_));
 sky130_fd_sc_hd__o211a_1 _11196_ (.A1(_04951_),
    .A2(_04952_),
    .B1(_04868_),
    .C1(_04870_),
    .X(_04955_));
 sky130_fd_sc_hd__a211oi_1 _11197_ (.A1(_04874_),
    .A2(_04878_),
    .B1(_04954_),
    .C1(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__o211a_1 _11198_ (.A1(_04954_),
    .A2(_04955_),
    .B1(_04874_),
    .C1(_04878_),
    .X(_04957_));
 sky130_fd_sc_hd__a211oi_1 _11199_ (.A1(_04838_),
    .A2(_04841_),
    .B1(_04956_),
    .C1(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__o211a_1 _11200_ (.A1(_04956_),
    .A2(_04957_),
    .B1(_04838_),
    .C1(_04841_),
    .X(_04959_));
 sky130_fd_sc_hd__o211a_1 _11201_ (.A1(_04958_),
    .A2(_04959_),
    .B1(_04880_),
    .C1(_04884_),
    .X(_04960_));
 sky130_fd_sc_hd__a211oi_1 _11202_ (.A1(_04880_),
    .A2(_04884_),
    .B1(_04958_),
    .C1(_04959_),
    .Y(_04961_));
 sky130_fd_sc_hd__nor2_1 _11203_ (.A(_04960_),
    .B(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__a21oi_1 _11204_ (.A1(_04889_),
    .A2(_04892_),
    .B1(_04887_),
    .Y(_04963_));
 sky130_fd_sc_hd__xnor2_1 _11205_ (.A(_04962_),
    .B(_04963_),
    .Y(net115));
 sky130_fd_sc_hd__nor2_4 _11206_ (.A(_04114_),
    .B(_04894_),
    .Y(_04965_));
 sky130_fd_sc_hd__a21oi_4 _11207_ (.A1(_04116_),
    .A2(_04894_),
    .B1(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__inv_2 _11208_ (.A(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__nand2b_1 _11209_ (.A_N(_04940_),
    .B(_04943_),
    .Y(_04968_));
 sky130_fd_sc_hd__o21bai_4 _11210_ (.A1(_04810_),
    .A2(_04893_),
    .B1_N(_04809_),
    .Y(_04969_));
 sky130_fd_sc_hd__and4_1 _11211_ (.A(net52),
    .B(net21),
    .C(net53),
    .D(net22),
    .X(_04970_));
 sky130_fd_sc_hd__a22o_1 _11212_ (.A1(net21),
    .A2(net53),
    .B1(net22),
    .B2(net52),
    .X(_04971_));
 sky130_fd_sc_hd__and2b_1 _11213_ (.A_N(_04970_),
    .B(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__nand2_1 _11214_ (.A(net20),
    .B(net54),
    .Y(_04973_));
 sky130_fd_sc_hd__xnor2_1 _11215_ (.A(_04972_),
    .B(_04973_),
    .Y(_04975_));
 sky130_fd_sc_hd__o21ba_1 _11216_ (.A1(_04902_),
    .A2(_04904_),
    .B1_N(_04901_),
    .X(_04976_));
 sky130_fd_sc_hd__nand2b_1 _11217_ (.A_N(_04976_),
    .B(_04975_),
    .Y(_04977_));
 sky130_fd_sc_hd__xnor2_1 _11218_ (.A(_04975_),
    .B(_04976_),
    .Y(_04978_));
 sky130_fd_sc_hd__and4b_1 _11219_ (.A_N(net18),
    .B(net19),
    .C(net56),
    .D(net57),
    .X(_04979_));
 sky130_fd_sc_hd__o2bb2a_1 _11220_ (.A1_N(net19),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net18),
    .X(_04980_));
 sky130_fd_sc_hd__nor2_1 _11221_ (.A(_04979_),
    .B(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__or2_1 _11222_ (.A(_04978_),
    .B(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__nand2_1 _11223_ (.A(_04978_),
    .B(_04981_),
    .Y(_04983_));
 sky130_fd_sc_hd__nand2_1 _11224_ (.A(_04982_),
    .B(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__and3_1 _11225_ (.A(_04907_),
    .B(_04915_),
    .C(_04984_),
    .X(_04986_));
 sky130_fd_sc_hd__a21oi_1 _11226_ (.A1(_04907_),
    .A2(_04915_),
    .B1(_04984_),
    .Y(_04987_));
 sky130_fd_sc_hd__or2_1 _11227_ (.A(_04986_),
    .B(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__and2_1 _11228_ (.A(_04911_),
    .B(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__nor2_1 _11229_ (.A(_04911_),
    .B(_04988_),
    .Y(_04990_));
 sky130_fd_sc_hd__or2_1 _11230_ (.A(_04989_),
    .B(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__a21o_1 _11231_ (.A1(_04924_),
    .A2(_04934_),
    .B1(_04933_),
    .X(_04992_));
 sky130_fd_sc_hd__and3_1 _11232_ (.A(net49),
    .B(net50),
    .C(net25),
    .X(_04993_));
 sky130_fd_sc_hd__o21ai_1 _11233_ (.A1(net49),
    .A2(net50),
    .B1(net25),
    .Y(_04994_));
 sky130_fd_sc_hd__nor2_2 _11234_ (.A(_04993_),
    .B(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__nand2_1 _11235_ (.A(net51),
    .B(net24),
    .Y(_04997_));
 sky130_fd_sc_hd__xor2_1 _11236_ (.A(_04995_),
    .B(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__xor2_1 _11237_ (.A(_04925_),
    .B(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__o21a_1 _11238_ (.A1(_04926_),
    .A2(_04930_),
    .B1(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__nor3_1 _11239_ (.A(_04926_),
    .B(_04930_),
    .C(_04999_),
    .Y(_05001_));
 sky130_fd_sc_hd__or2_1 _11240_ (.A(_05000_),
    .B(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__nor2_1 _11241_ (.A(_04923_),
    .B(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__xor2_1 _11242_ (.A(_04923_),
    .B(_05002_),
    .X(_05004_));
 sky130_fd_sc_hd__xnor2_1 _11243_ (.A(_04992_),
    .B(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__a21oi_1 _11244_ (.A1(_04936_),
    .A2(_04938_),
    .B1(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__and3_1 _11245_ (.A(_04936_),
    .B(_04938_),
    .C(_05005_),
    .X(_05008_));
 sky130_fd_sc_hd__or2_1 _11246_ (.A(_05006_),
    .B(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__xnor2_1 _11247_ (.A(_04991_),
    .B(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__and2b_1 _11248_ (.A_N(_05010_),
    .B(_04969_),
    .X(_05011_));
 sky130_fd_sc_hd__xor2_1 _11249_ (.A(_04969_),
    .B(_05010_),
    .X(_05012_));
 sky130_fd_sc_hd__and2b_1 _11250_ (.A_N(_05012_),
    .B(_04968_),
    .X(_05013_));
 sky130_fd_sc_hd__xor2_1 _11251_ (.A(_04968_),
    .B(_05012_),
    .X(_05014_));
 sky130_fd_sc_hd__xnor2_1 _11252_ (.A(_04966_),
    .B(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__or2_1 _11253_ (.A(_04896_),
    .B(_04950_),
    .X(_05016_));
 sky130_fd_sc_hd__nand2_1 _11254_ (.A(_05015_),
    .B(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__or2_1 _11255_ (.A(_05015_),
    .B(_05016_),
    .X(_05019_));
 sky130_fd_sc_hd__nand2_1 _11256_ (.A(_05017_),
    .B(_05019_),
    .Y(_05020_));
 sky130_fd_sc_hd__nand2_1 _11257_ (.A(_04945_),
    .B(_04947_),
    .Y(_05021_));
 sky130_fd_sc_hd__nand2b_1 _11258_ (.A_N(_05020_),
    .B(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__nand2b_1 _11259_ (.A_N(_05021_),
    .B(_05020_),
    .Y(_05023_));
 sky130_fd_sc_hd__o211a_1 _11260_ (.A1(_04951_),
    .A2(_04954_),
    .B1(_05022_),
    .C1(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__a211oi_1 _11261_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_04951_),
    .C1(_04954_),
    .Y(_05025_));
 sky130_fd_sc_hd__or2_1 _11262_ (.A(_05024_),
    .B(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__o21ba_1 _11263_ (.A1(_04830_),
    .A2(_04919_),
    .B1_N(_04918_),
    .X(_05027_));
 sky130_fd_sc_hd__xnor2_1 _11264_ (.A(_05026_),
    .B(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__or2_1 _11265_ (.A(_04956_),
    .B(_04958_),
    .X(_05030_));
 sky130_fd_sc_hd__and2b_1 _11266_ (.A_N(_05028_),
    .B(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__xnor2_1 _11267_ (.A(_05028_),
    .B(_05030_),
    .Y(_05032_));
 sky130_fd_sc_hd__nand2_1 _11268_ (.A(_04889_),
    .B(_04962_),
    .Y(_05033_));
 sky130_fd_sc_hd__nor2_1 _11269_ (.A(_04891_),
    .B(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__nand2_1 _11270_ (.A(_04714_),
    .B(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__a211o_1 _11271_ (.A1(_03350_),
    .A2(_04339_),
    .B1(_05035_),
    .C1(_04338_),
    .X(_05036_));
 sky130_fd_sc_hd__nand2_1 _11272_ (.A(_04713_),
    .B(_05034_),
    .Y(_05037_));
 sky130_fd_sc_hd__o21bai_1 _11273_ (.A1(_04887_),
    .A2(_04961_),
    .B1_N(_04960_),
    .Y(_05038_));
 sky130_fd_sc_hd__o211a_1 _11274_ (.A1(_04890_),
    .A2(_05033_),
    .B1(_05037_),
    .C1(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__nand2_1 _11275_ (.A(_05036_),
    .B(_05039_),
    .Y(_05041_));
 sky130_fd_sc_hd__xor2_1 _11276_ (.A(_05032_),
    .B(_05041_),
    .X(net116));
 sky130_fd_sc_hd__o21bai_1 _11277_ (.A1(_04991_),
    .A2(_05008_),
    .B1_N(_05006_),
    .Y(_05042_));
 sky130_fd_sc_hd__and4_1 _11278_ (.A(net52),
    .B(net53),
    .C(net22),
    .D(net24),
    .X(_05043_));
 sky130_fd_sc_hd__a22oi_1 _11279_ (.A1(net53),
    .A2(net22),
    .B1(net24),
    .B2(net52),
    .Y(_05044_));
 sky130_fd_sc_hd__nor2_1 _11280_ (.A(_05043_),
    .B(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand2_1 _11281_ (.A(net21),
    .B(net54),
    .Y(_05046_));
 sky130_fd_sc_hd__xnor2_1 _11282_ (.A(_05045_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__a31o_1 _11283_ (.A1(net20),
    .A2(net54),
    .A3(_04971_),
    .B1(_04970_),
    .X(_05048_));
 sky130_fd_sc_hd__nor2_1 _11284_ (.A(_05047_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__and2_1 _11285_ (.A(_05047_),
    .B(_05048_),
    .X(_05051_));
 sky130_fd_sc_hd__nor2_1 _11286_ (.A(_05049_),
    .B(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__and4b_1 _11287_ (.A_N(net19),
    .B(net20),
    .C(net56),
    .D(net57),
    .X(_05053_));
 sky130_fd_sc_hd__o2bb2a_1 _11288_ (.A1_N(net20),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net19),
    .X(_05054_));
 sky130_fd_sc_hd__nor2_1 _11289_ (.A(_05053_),
    .B(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__xnor2_1 _11290_ (.A(_05052_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__and3_1 _11291_ (.A(_04977_),
    .B(_04983_),
    .C(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__a21o_1 _11292_ (.A1(_04977_),
    .A2(_04983_),
    .B1(_05056_),
    .X(_05058_));
 sky130_fd_sc_hd__and2b_1 _11293_ (.A_N(_05057_),
    .B(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__or2_1 _11294_ (.A(_04979_),
    .B(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__nand2_1 _11295_ (.A(_04979_),
    .B(_05059_),
    .Y(_05062_));
 sky130_fd_sc_hd__nand2_1 _11296_ (.A(_05060_),
    .B(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__o21ba_1 _11297_ (.A1(_04925_),
    .A2(_04998_),
    .B1_N(_05000_),
    .X(_05064_));
 sky130_fd_sc_hd__a31o_1 _11298_ (.A1(net51),
    .A2(net24),
    .A3(_04995_),
    .B1(_04993_),
    .X(_05065_));
 sky130_fd_sc_hd__a21oi_1 _11299_ (.A1(net51),
    .A2(net25),
    .B1(_04995_),
    .Y(_05066_));
 sky130_fd_sc_hd__a21o_1 _11300_ (.A1(net51),
    .A2(_04995_),
    .B1(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__or2_1 _11301_ (.A(_04925_),
    .B(_05067_),
    .X(_05068_));
 sky130_fd_sc_hd__xnor2_1 _11302_ (.A(_04925_),
    .B(_05067_),
    .Y(_05069_));
 sky130_fd_sc_hd__nand2b_1 _11303_ (.A_N(_05069_),
    .B(_05065_),
    .Y(_05070_));
 sky130_fd_sc_hd__xor2_1 _11304_ (.A(_05065_),
    .B(_05069_),
    .X(_05071_));
 sky130_fd_sc_hd__or2_1 _11305_ (.A(_04923_),
    .B(_05071_),
    .X(_05073_));
 sky130_fd_sc_hd__xor2_1 _11306_ (.A(_04923_),
    .B(_05071_),
    .X(_05074_));
 sky130_fd_sc_hd__nand2b_1 _11307_ (.A_N(_05064_),
    .B(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__xnor2_1 _11308_ (.A(_05064_),
    .B(_05074_),
    .Y(_05076_));
 sky130_fd_sc_hd__a21o_1 _11309_ (.A1(_04992_),
    .A2(_05004_),
    .B1(_05003_),
    .X(_05077_));
 sky130_fd_sc_hd__xnor2_1 _11310_ (.A(_05076_),
    .B(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__or2_1 _11311_ (.A(_05063_),
    .B(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__xnor2_1 _11312_ (.A(_05063_),
    .B(_05078_),
    .Y(_05080_));
 sky130_fd_sc_hd__and2b_1 _11313_ (.A_N(_05080_),
    .B(_04969_),
    .X(_05081_));
 sky130_fd_sc_hd__xor2_1 _11314_ (.A(_04969_),
    .B(_05080_),
    .X(_05082_));
 sky130_fd_sc_hd__and2b_1 _11315_ (.A_N(_05082_),
    .B(_05042_),
    .X(_05084_));
 sky130_fd_sc_hd__xor2_1 _11316_ (.A(_05042_),
    .B(_05082_),
    .X(_05085_));
 sky130_fd_sc_hd__xnor2_1 _11317_ (.A(_04966_),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__o21bai_1 _11318_ (.A1(_04967_),
    .A2(_05014_),
    .B1_N(_04965_),
    .Y(_05087_));
 sky130_fd_sc_hd__nand2_1 _11319_ (.A(_05086_),
    .B(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__or2_1 _11320_ (.A(_05086_),
    .B(_05087_),
    .X(_05089_));
 sky130_fd_sc_hd__and2_1 _11321_ (.A(_05088_),
    .B(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__o21a_1 _11322_ (.A1(_05011_),
    .A2(_05013_),
    .B1(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__o21ai_1 _11323_ (.A1(_05011_),
    .A2(_05013_),
    .B1(_05090_),
    .Y(_05092_));
 sky130_fd_sc_hd__nor3_1 _11324_ (.A(_05011_),
    .B(_05013_),
    .C(_05090_),
    .Y(_05093_));
 sky130_fd_sc_hd__a211o_1 _11325_ (.A1(_05017_),
    .A2(_05022_),
    .B1(_05091_),
    .C1(_05093_),
    .X(_05095_));
 sky130_fd_sc_hd__o211ai_2 _11326_ (.A1(_05091_),
    .A2(_05093_),
    .B1(_05017_),
    .C1(_05022_),
    .Y(_05096_));
 sky130_fd_sc_hd__o211ai_2 _11327_ (.A1(_04987_),
    .A2(_04990_),
    .B1(_05095_),
    .C1(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__a211o_1 _11328_ (.A1(_05095_),
    .A2(_05096_),
    .B1(_04987_),
    .C1(_04990_),
    .X(_05098_));
 sky130_fd_sc_hd__nand2_1 _11329_ (.A(_05097_),
    .B(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__o21bai_2 _11330_ (.A1(_05025_),
    .A2(_05027_),
    .B1_N(_05024_),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2b_1 _11331_ (.A_N(_05100_),
    .B(_05099_),
    .Y(_05101_));
 sky130_fd_sc_hd__xnor2_1 _11332_ (.A(_05099_),
    .B(_05100_),
    .Y(_05102_));
 sky130_fd_sc_hd__a21oi_1 _11333_ (.A1(_05032_),
    .A2(_05041_),
    .B1(_05031_),
    .Y(_05103_));
 sky130_fd_sc_hd__xnor2_1 _11334_ (.A(_05102_),
    .B(_05103_),
    .Y(net117));
 sky130_fd_sc_hd__a21bo_1 _11335_ (.A1(_05076_),
    .A2(_05077_),
    .B1_N(_05079_),
    .X(_05105_));
 sky130_fd_sc_hd__and3_1 _11336_ (.A(net52),
    .B(net53),
    .C(net25),
    .X(_05106_));
 sky130_fd_sc_hd__and2_1 _11337_ (.A(net24),
    .B(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__a22oi_1 _11338_ (.A1(net53),
    .A2(net24),
    .B1(net25),
    .B2(net52),
    .Y(_05108_));
 sky130_fd_sc_hd__nor2_1 _11339_ (.A(_05107_),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__a21oi_1 _11340_ (.A1(net22),
    .A2(net54),
    .B1(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hd__and3_1 _11341_ (.A(net22),
    .B(net54),
    .C(_05109_),
    .X(_05111_));
 sky130_fd_sc_hd__or2_1 _11342_ (.A(_05110_),
    .B(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__o21ba_1 _11343_ (.A1(_05044_),
    .A2(_05046_),
    .B1_N(_05043_),
    .X(_05113_));
 sky130_fd_sc_hd__xnor2_1 _11344_ (.A(_05112_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__and4b_1 _11345_ (.A_N(net20),
    .B(net21),
    .C(net56),
    .D(net57),
    .X(_05116_));
 sky130_fd_sc_hd__o2bb2a_1 _11346_ (.A1_N(net21),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net20),
    .X(_05117_));
 sky130_fd_sc_hd__nor2_1 _11347_ (.A(_05116_),
    .B(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__xnor2_1 _11348_ (.A(_05114_),
    .B(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__a21oi_1 _11349_ (.A1(_05052_),
    .A2(_05055_),
    .B1(_05051_),
    .Y(_05120_));
 sky130_fd_sc_hd__nand2b_1 _11350_ (.A_N(_05120_),
    .B(_05119_),
    .Y(_05121_));
 sky130_fd_sc_hd__xnor2_1 _11351_ (.A(_05119_),
    .B(_05120_),
    .Y(_05122_));
 sky130_fd_sc_hd__or2_1 _11352_ (.A(_05053_),
    .B(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__nand2_1 _11353_ (.A(_05053_),
    .B(_05122_),
    .Y(_05124_));
 sky130_fd_sc_hd__nand2_1 _11354_ (.A(_05123_),
    .B(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__nand2_1 _11355_ (.A(_05068_),
    .B(_05070_),
    .Y(_05127_));
 sky130_fd_sc_hd__a21oi_2 _11356_ (.A1(net51),
    .A2(_04995_),
    .B1(_04993_),
    .Y(_05128_));
 sky130_fd_sc_hd__xor2_1 _11357_ (.A(_05069_),
    .B(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__xnor2_1 _11358_ (.A(_04923_),
    .B(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__xnor2_1 _11359_ (.A(_05127_),
    .B(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__a21oi_2 _11360_ (.A1(_05073_),
    .A2(_05075_),
    .B1(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__and3_1 _11361_ (.A(_05073_),
    .B(_05075_),
    .C(_05131_),
    .X(_05133_));
 sky130_fd_sc_hd__or3_1 _11362_ (.A(_05125_),
    .B(_05132_),
    .C(_05133_),
    .X(_05134_));
 sky130_fd_sc_hd__inv_2 _11363_ (.A(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__o21ai_1 _11364_ (.A1(_05132_),
    .A2(_05133_),
    .B1(_05125_),
    .Y(_05136_));
 sky130_fd_sc_hd__and3_1 _11365_ (.A(_04969_),
    .B(_05134_),
    .C(_05136_),
    .X(_05138_));
 sky130_fd_sc_hd__a21oi_1 _11366_ (.A1(_05134_),
    .A2(_05136_),
    .B1(_04969_),
    .Y(_05139_));
 sky130_fd_sc_hd__or2_1 _11367_ (.A(_05138_),
    .B(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__and2b_1 _11368_ (.A_N(_05140_),
    .B(_05105_),
    .X(_05141_));
 sky130_fd_sc_hd__xor2_1 _11369_ (.A(_05105_),
    .B(_05140_),
    .X(_05142_));
 sky130_fd_sc_hd__xnor2_1 _11370_ (.A(_04966_),
    .B(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__o21bai_1 _11371_ (.A1(_04967_),
    .A2(_05085_),
    .B1_N(_04965_),
    .Y(_05144_));
 sky130_fd_sc_hd__nand2_1 _11372_ (.A(_05143_),
    .B(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__or2_1 _11373_ (.A(_05143_),
    .B(_05144_),
    .X(_05146_));
 sky130_fd_sc_hd__and2_1 _11374_ (.A(_05145_),
    .B(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__o21ai_2 _11375_ (.A1(_05081_),
    .A2(_05084_),
    .B1(_05147_),
    .Y(_05149_));
 sky130_fd_sc_hd__or3_1 _11376_ (.A(_05081_),
    .B(_05084_),
    .C(_05147_),
    .X(_05150_));
 sky130_fd_sc_hd__nand2_1 _11377_ (.A(_05149_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__a21oi_2 _11378_ (.A1(_05088_),
    .A2(_05092_),
    .B1(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__and3_1 _11379_ (.A(_05088_),
    .B(_05092_),
    .C(_05151_),
    .X(_05153_));
 sky130_fd_sc_hd__a211oi_2 _11380_ (.A1(_05058_),
    .A2(_05062_),
    .B1(_05152_),
    .C1(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__o211a_1 _11381_ (.A1(_05152_),
    .A2(_05153_),
    .B1(_05058_),
    .C1(_05062_),
    .X(_05155_));
 sky130_fd_sc_hd__a211oi_1 _11382_ (.A1(_05095_),
    .A2(_05097_),
    .B1(_05154_),
    .C1(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__o211ai_1 _11383_ (.A1(_05154_),
    .A2(_05155_),
    .B1(_05095_),
    .C1(_05097_),
    .Y(_05157_));
 sky130_fd_sc_hd__nand2b_1 _11384_ (.A_N(_05156_),
    .B(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__nand2_1 _11385_ (.A(_05032_),
    .B(_05102_),
    .Y(_05160_));
 sky130_fd_sc_hd__a21oi_2 _11386_ (.A1(_05036_),
    .A2(_05039_),
    .B1(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__and2_1 _11387_ (.A(_05031_),
    .B(_05101_),
    .X(_05162_));
 sky130_fd_sc_hd__a31o_1 _11388_ (.A1(_05097_),
    .A2(_05098_),
    .A3(_05100_),
    .B1(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__nor2_1 _11389_ (.A(_05161_),
    .B(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__xor2_1 _11390_ (.A(_05158_),
    .B(_05164_),
    .X(net118));
 sky130_fd_sc_hd__o21ai_1 _11391_ (.A1(net52),
    .A2(net53),
    .B1(net25),
    .Y(_05165_));
 sky130_fd_sc_hd__nor2_1 _11392_ (.A(_05106_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__nand2_1 _11393_ (.A(net54),
    .B(net24),
    .Y(_05167_));
 sky130_fd_sc_hd__xnor2_1 _11394_ (.A(_05166_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__or3_1 _11395_ (.A(_05107_),
    .B(_05111_),
    .C(_05168_),
    .X(_05170_));
 sky130_fd_sc_hd__o21ai_1 _11396_ (.A1(_05107_),
    .A2(_05111_),
    .B1(_05168_),
    .Y(_05171_));
 sky130_fd_sc_hd__nand2_1 _11397_ (.A(_05170_),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__and4b_1 _11398_ (.A_N(net21),
    .B(net22),
    .C(net56),
    .D(net57),
    .X(_05173_));
 sky130_fd_sc_hd__inv_2 _11399_ (.A(_05173_),
    .Y(_05174_));
 sky130_fd_sc_hd__o2bb2a_1 _11400_ (.A1_N(net22),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net21),
    .X(_05175_));
 sky130_fd_sc_hd__o21ai_1 _11401_ (.A1(_05173_),
    .A2(_05175_),
    .B1(_05172_),
    .Y(_05176_));
 sky130_fd_sc_hd__or3_1 _11402_ (.A(_05172_),
    .B(_05173_),
    .C(_05175_),
    .X(_05177_));
 sky130_fd_sc_hd__and2_1 _11403_ (.A(_05176_),
    .B(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__o32a_1 _11404_ (.A1(_05114_),
    .A2(_05116_),
    .A3(_05117_),
    .B1(_05113_),
    .B2(_05112_),
    .X(_05179_));
 sky130_fd_sc_hd__and2b_1 _11405_ (.A_N(_05179_),
    .B(_05178_),
    .X(_05181_));
 sky130_fd_sc_hd__xnor2_1 _11406_ (.A(_05178_),
    .B(_05179_),
    .Y(_05182_));
 sky130_fd_sc_hd__xnor2_1 _11407_ (.A(_05116_),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__and4_2 _11408_ (.A(_04923_),
    .B(_04925_),
    .C(_05067_),
    .D(_05128_),
    .X(_05184_));
 sky130_fd_sc_hd__nor2_1 _11409_ (.A(_05132_),
    .B(_05184_),
    .Y(_05185_));
 sky130_fd_sc_hd__xnor2_1 _11410_ (.A(_05183_),
    .B(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__xor2_1 _11411_ (.A(_04969_),
    .B(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__o21a_1 _11412_ (.A1(_05132_),
    .A2(_05135_),
    .B1(_05187_),
    .X(_05188_));
 sky130_fd_sc_hd__nor3_1 _11413_ (.A(_05132_),
    .B(_05135_),
    .C(_05187_),
    .Y(_05189_));
 sky130_fd_sc_hd__nor2_1 _11414_ (.A(_05188_),
    .B(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__xnor2_1 _11415_ (.A(_04966_),
    .B(_05190_),
    .Y(_05192_));
 sky130_fd_sc_hd__o21bai_1 _11416_ (.A1(_04967_),
    .A2(_05142_),
    .B1_N(_04965_),
    .Y(_05193_));
 sky130_fd_sc_hd__and2b_1 _11417_ (.A_N(_05192_),
    .B(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__xnor2_1 _11418_ (.A(_05192_),
    .B(_05193_),
    .Y(_05195_));
 sky130_fd_sc_hd__o21a_1 _11419_ (.A1(_05138_),
    .A2(_05141_),
    .B1(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__nor3_1 _11420_ (.A(_05138_),
    .B(_05141_),
    .C(_05195_),
    .Y(_05197_));
 sky130_fd_sc_hd__a211oi_2 _11421_ (.A1(_05145_),
    .A2(_05149_),
    .B1(_05196_),
    .C1(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__o211a_1 _11422_ (.A1(_05196_),
    .A2(_05197_),
    .B1(_05145_),
    .C1(_05149_),
    .X(_05199_));
 sky130_fd_sc_hd__a211oi_2 _11423_ (.A1(_05121_),
    .A2(_05124_),
    .B1(_05198_),
    .C1(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__inv_2 _11424_ (.A(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__o211ai_1 _11425_ (.A1(_05198_),
    .A2(_05199_),
    .B1(_05121_),
    .C1(_05124_),
    .Y(_05203_));
 sky130_fd_sc_hd__a211o_1 _11426_ (.A1(_05201_),
    .A2(_05203_),
    .B1(_05152_),
    .C1(_05154_),
    .X(_05204_));
 sky130_fd_sc_hd__inv_2 _11427_ (.A(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__o211a_1 _11428_ (.A1(_05152_),
    .A2(_05154_),
    .B1(_05201_),
    .C1(_05203_),
    .X(_05206_));
 sky130_fd_sc_hd__nor2_1 _11429_ (.A(_05205_),
    .B(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__o21ba_1 _11430_ (.A1(_05158_),
    .A2(_05164_),
    .B1_N(_05156_),
    .X(_05208_));
 sky130_fd_sc_hd__xnor2_1 _11431_ (.A(_05207_),
    .B(_05208_),
    .Y(net119));
 sky130_fd_sc_hd__nor3_1 _11432_ (.A(_04923_),
    .B(_05068_),
    .C(_05128_),
    .Y(_05209_));
 sky130_fd_sc_hd__or3_1 _11433_ (.A(_04923_),
    .B(_05068_),
    .C(_05128_),
    .X(_05210_));
 sky130_fd_sc_hd__o31ai_1 _11434_ (.A1(_05132_),
    .A2(_05183_),
    .A3(_05184_),
    .B1(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__and4b_1 _11435_ (.A_N(net22),
    .B(net24),
    .C(net56),
    .D(net57),
    .X(_05213_));
 sky130_fd_sc_hd__o2bb2a_1 _11436_ (.A1_N(net24),
    .A2_N(net56),
    .B1(_00287_),
    .B2(net22),
    .X(_05214_));
 sky130_fd_sc_hd__nor2_1 _11437_ (.A(_05213_),
    .B(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__nand2_1 _11438_ (.A(net54),
    .B(net25),
    .Y(_05216_));
 sky130_fd_sc_hd__xnor2_1 _11439_ (.A(_05166_),
    .B(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__and2_1 _11440_ (.A(net54),
    .B(_05106_),
    .X(_05218_));
 sky130_fd_sc_hd__nand2_1 _11441_ (.A(net54),
    .B(_05106_),
    .Y(_05219_));
 sky130_fd_sc_hd__a311o_1 _11442_ (.A1(net54),
    .A2(net24),
    .A3(_05166_),
    .B1(_05217_),
    .C1(_05106_),
    .X(_05220_));
 sky130_fd_sc_hd__and2_1 _11443_ (.A(_05219_),
    .B(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__xnor2_1 _11444_ (.A(_05215_),
    .B(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__nand3_1 _11445_ (.A(_05171_),
    .B(_05177_),
    .C(_05222_),
    .Y(_05224_));
 sky130_fd_sc_hd__a21o_1 _11446_ (.A1(_05171_),
    .A2(_05177_),
    .B1(_05222_),
    .X(_05225_));
 sky130_fd_sc_hd__nand2_1 _11447_ (.A(_05224_),
    .B(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__xnor2_1 _11448_ (.A(_05174_),
    .B(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__nor2_2 _11449_ (.A(_05184_),
    .B(_05209_),
    .Y(_05228_));
 sky130_fd_sc_hd__or3_1 _11450_ (.A(_05184_),
    .B(_05209_),
    .C(_05227_),
    .X(_05229_));
 sky130_fd_sc_hd__xnor2_1 _11451_ (.A(_05227_),
    .B(_05228_),
    .Y(_05230_));
 sky130_fd_sc_hd__xnor2_1 _11452_ (.A(_04969_),
    .B(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__and2b_1 _11453_ (.A_N(_05231_),
    .B(_05211_),
    .X(_05232_));
 sky130_fd_sc_hd__xnor2_1 _11454_ (.A(_05211_),
    .B(_05231_),
    .Y(_05233_));
 sky130_fd_sc_hd__xnor2_1 _11455_ (.A(_04967_),
    .B(_05233_),
    .Y(_05235_));
 sky130_fd_sc_hd__a21o_1 _11456_ (.A1(_04966_),
    .A2(_05190_),
    .B1(_04965_),
    .X(_05236_));
 sky130_fd_sc_hd__nand2_1 _11457_ (.A(_05235_),
    .B(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__or2_1 _11458_ (.A(_05235_),
    .B(_05236_),
    .X(_05238_));
 sky130_fd_sc_hd__and2_1 _11459_ (.A(_05237_),
    .B(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__a21oi_1 _11460_ (.A1(_04969_),
    .A2(_05186_),
    .B1(_05188_),
    .Y(_05240_));
 sky130_fd_sc_hd__nand2b_1 _11461_ (.A_N(_05240_),
    .B(_05239_),
    .Y(_05241_));
 sky130_fd_sc_hd__xnor2_1 _11462_ (.A(_05239_),
    .B(_05240_),
    .Y(_05242_));
 sky130_fd_sc_hd__nor2_1 _11463_ (.A(_05194_),
    .B(_05196_),
    .Y(_05243_));
 sky130_fd_sc_hd__and2b_1 _11464_ (.A_N(_05243_),
    .B(_05242_),
    .X(_05244_));
 sky130_fd_sc_hd__xnor2_1 _11465_ (.A(_05242_),
    .B(_05243_),
    .Y(_05246_));
 sky130_fd_sc_hd__a21oi_1 _11466_ (.A1(_05116_),
    .A2(_05182_),
    .B1(_05181_),
    .Y(_05247_));
 sky130_fd_sc_hd__and2b_1 _11467_ (.A_N(_05247_),
    .B(_05246_),
    .X(_05248_));
 sky130_fd_sc_hd__xnor2_1 _11468_ (.A(_05246_),
    .B(_05247_),
    .Y(_05249_));
 sky130_fd_sc_hd__o21ai_1 _11469_ (.A1(_05198_),
    .A2(_05200_),
    .B1(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__or3_1 _11470_ (.A(_05198_),
    .B(_05200_),
    .C(_05249_),
    .X(_05251_));
 sky130_fd_sc_hd__nand2_1 _11471_ (.A(_05250_),
    .B(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hd__inv_2 _11472_ (.A(_05252_),
    .Y(_05253_));
 sky130_fd_sc_hd__a21o_1 _11473_ (.A1(_05156_),
    .A2(_05204_),
    .B1(_05206_),
    .X(_05254_));
 sky130_fd_sc_hd__a21o_1 _11474_ (.A1(_05157_),
    .A2(_05204_),
    .B1(_05206_),
    .X(_05255_));
 sky130_fd_sc_hd__o31a_1 _11475_ (.A1(_05161_),
    .A2(_05163_),
    .A3(_05254_),
    .B1(_05255_),
    .X(_05257_));
 sky130_fd_sc_hd__o311ai_2 _11476_ (.A1(_05161_),
    .A2(_05163_),
    .A3(_05254_),
    .B1(_05255_),
    .C1(_05253_),
    .Y(_05258_));
 sky130_fd_sc_hd__or2_1 _11477_ (.A(_05253_),
    .B(_05257_),
    .X(_05259_));
 sky130_fd_sc_hd__and2_1 _11478_ (.A(_05258_),
    .B(_05259_),
    .X(net121));
 sky130_fd_sc_hd__nand2_1 _11479_ (.A(_05165_),
    .B(_05216_),
    .Y(_05260_));
 sky130_fd_sc_hd__nand2_1 _11480_ (.A(_05219_),
    .B(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__o2bb2a_1 _11481_ (.A1_N(net56),
    .A2_N(net25),
    .B1(_00287_),
    .B2(net24),
    .X(_05262_));
 sky130_fd_sc_hd__and4b_1 _11482_ (.A_N(net24),
    .B(net56),
    .C(net57),
    .D(net25),
    .X(_05263_));
 sky130_fd_sc_hd__o21ai_1 _11483_ (.A1(_05262_),
    .A2(_05263_),
    .B1(_05261_),
    .Y(_05264_));
 sky130_fd_sc_hd__or3_1 _11484_ (.A(_05261_),
    .B(_05262_),
    .C(_05263_),
    .X(_05265_));
 sky130_fd_sc_hd__and2_1 _11485_ (.A(_05264_),
    .B(_05265_),
    .X(_05267_));
 sky130_fd_sc_hd__a21o_1 _11486_ (.A1(_05215_),
    .A2(_05220_),
    .B1(_05218_),
    .X(_05268_));
 sky130_fd_sc_hd__nor2_1 _11487_ (.A(_05267_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__and2_1 _11488_ (.A(_05267_),
    .B(_05268_),
    .X(_05270_));
 sky130_fd_sc_hd__nor2_1 _11489_ (.A(_05269_),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__xnor2_1 _11490_ (.A(_05213_),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__xor2_1 _11491_ (.A(_05228_),
    .B(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__inv_2 _11492_ (.A(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__xor2_1 _11493_ (.A(_04969_),
    .B(_05273_),
    .X(_05275_));
 sky130_fd_sc_hd__a21oi_1 _11494_ (.A1(_05210_),
    .A2(_05229_),
    .B1(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__and3_1 _11495_ (.A(_05210_),
    .B(_05229_),
    .C(_05275_),
    .X(_05278_));
 sky130_fd_sc_hd__or2_1 _11496_ (.A(_05276_),
    .B(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__and2_1 _11497_ (.A(_04967_),
    .B(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__nor2_1 _11498_ (.A(_04967_),
    .B(_05279_),
    .Y(_05281_));
 sky130_fd_sc_hd__or2_1 _11499_ (.A(_05280_),
    .B(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__a21o_1 _11500_ (.A1(_04966_),
    .A2(_05233_),
    .B1(_04965_),
    .X(_05283_));
 sky130_fd_sc_hd__nand2b_1 _11501_ (.A_N(_05282_),
    .B(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__nand2b_1 _11502_ (.A_N(_05283_),
    .B(_05282_),
    .Y(_05285_));
 sky130_fd_sc_hd__nand2_1 _11503_ (.A(_05284_),
    .B(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__a21oi_1 _11504_ (.A1(_04969_),
    .A2(_05230_),
    .B1(_05232_),
    .Y(_05287_));
 sky130_fd_sc_hd__xnor2_1 _11505_ (.A(_05286_),
    .B(_05287_),
    .Y(_05289_));
 sky130_fd_sc_hd__a21oi_1 _11506_ (.A1(_05237_),
    .A2(_05241_),
    .B1(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__and3_1 _11507_ (.A(_05237_),
    .B(_05241_),
    .C(_05289_),
    .X(_05291_));
 sky130_fd_sc_hd__or2_1 _11508_ (.A(_05290_),
    .B(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__o21ai_1 _11509_ (.A1(_05174_),
    .A2(_05226_),
    .B1(_05225_),
    .Y(_05293_));
 sky130_fd_sc_hd__and2b_1 _11510_ (.A_N(_05292_),
    .B(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__xnor2_1 _11511_ (.A(_05292_),
    .B(_05293_),
    .Y(_05295_));
 sky130_fd_sc_hd__o21ai_1 _11512_ (.A1(_05244_),
    .A2(_05248_),
    .B1(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__nor3_1 _11513_ (.A(_05244_),
    .B(_05248_),
    .C(_05295_),
    .Y(_05297_));
 sky130_fd_sc_hd__inv_2 _11514_ (.A(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__nand2_1 _11515_ (.A(_05296_),
    .B(_05298_),
    .Y(_05300_));
 sky130_fd_sc_hd__nand2_1 _11516_ (.A(_05250_),
    .B(_05258_),
    .Y(_05301_));
 sky130_fd_sc_hd__xnor2_1 _11517_ (.A(_05300_),
    .B(_05301_),
    .Y(net122));
 sky130_fd_sc_hd__o21ai_1 _11518_ (.A1(_05184_),
    .A2(_05272_),
    .B1(_05210_),
    .Y(_05302_));
 sky130_fd_sc_hd__mux2_1 _11519_ (.A0(net57),
    .A1(net56),
    .S(net25),
    .X(_05303_));
 sky130_fd_sc_hd__xor2_1 _11520_ (.A(_05261_),
    .B(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__a21oi_1 _11521_ (.A1(_05219_),
    .A2(_05265_),
    .B1(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__and3_1 _11522_ (.A(_05219_),
    .B(_05265_),
    .C(_05304_),
    .X(_05306_));
 sky130_fd_sc_hd__or2_1 _11523_ (.A(_05305_),
    .B(_05306_),
    .X(_05307_));
 sky130_fd_sc_hd__inv_2 _11524_ (.A(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__xor2_1 _11525_ (.A(_05263_),
    .B(_05307_),
    .X(_05310_));
 sky130_fd_sc_hd__xnor2_1 _11526_ (.A(_05228_),
    .B(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__xnor2_1 _11527_ (.A(_05302_),
    .B(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__xor2_1 _11528_ (.A(_04969_),
    .B(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__xnor2_1 _11529_ (.A(_04966_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__o21ai_1 _11530_ (.A1(_04965_),
    .A2(_05281_),
    .B1(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__or3_1 _11531_ (.A(_04965_),
    .B(_05281_),
    .C(_05314_),
    .X(_05316_));
 sky130_fd_sc_hd__nand2_1 _11532_ (.A(_05315_),
    .B(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__a21oi_1 _11533_ (.A1(_04969_),
    .A2(_05274_),
    .B1(_05276_),
    .Y(_05318_));
 sky130_fd_sc_hd__xor2_1 _11534_ (.A(_05317_),
    .B(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__o21a_1 _11535_ (.A1(_05286_),
    .A2(_05287_),
    .B1(_05284_),
    .X(_05321_));
 sky130_fd_sc_hd__nand2b_1 _11536_ (.A_N(_05321_),
    .B(_05319_),
    .Y(_05322_));
 sky130_fd_sc_hd__nand2b_1 _11537_ (.A_N(_05319_),
    .B(_05321_),
    .Y(_05323_));
 sky130_fd_sc_hd__nand2_1 _11538_ (.A(_05322_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__a21oi_1 _11539_ (.A1(_05213_),
    .A2(_05271_),
    .B1(_05270_),
    .Y(_05325_));
 sky130_fd_sc_hd__xor2_1 _11540_ (.A(_05324_),
    .B(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__o21a_1 _11541_ (.A1(_05290_),
    .A2(_05294_),
    .B1(_05326_),
    .X(_05327_));
 sky130_fd_sc_hd__o21ai_1 _11542_ (.A1(_05290_),
    .A2(_05294_),
    .B1(_05326_),
    .Y(_05328_));
 sky130_fd_sc_hd__nor3_1 _11543_ (.A(_05290_),
    .B(_05294_),
    .C(_05326_),
    .Y(_05329_));
 sky130_fd_sc_hd__nor2_1 _11544_ (.A(_05327_),
    .B(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__a31o_1 _11545_ (.A1(_05250_),
    .A2(_05258_),
    .A3(_05296_),
    .B1(_05297_),
    .X(_05332_));
 sky130_fd_sc_hd__xnor2_1 _11546_ (.A(_05330_),
    .B(_05332_),
    .Y(net123));
 sky130_fd_sc_hd__o21ai_1 _11547_ (.A1(_05324_),
    .A2(_05325_),
    .B1(_05322_),
    .Y(_05333_));
 sky130_fd_sc_hd__o21a_1 _11548_ (.A1(_05317_),
    .A2(_05318_),
    .B1(_05315_),
    .X(_05334_));
 sky130_fd_sc_hd__a21o_1 _11549_ (.A1(_04966_),
    .A2(_05313_),
    .B1(_04965_),
    .X(_05335_));
 sky130_fd_sc_hd__mux2_1 _11550_ (.A0(_05311_),
    .A1(_04969_),
    .S(_05302_),
    .X(_05336_));
 sky130_fd_sc_hd__o21ba_1 _11551_ (.A1(_04969_),
    .A2(_05311_),
    .B1_N(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__a21o_1 _11552_ (.A1(_05228_),
    .A2(_05310_),
    .B1(_05209_),
    .X(_05338_));
 sky130_fd_sc_hd__or3_1 _11553_ (.A(_05218_),
    .B(_05260_),
    .C(_05303_),
    .X(_05339_));
 sky130_fd_sc_hd__a21oi_1 _11554_ (.A1(_05263_),
    .A2(_05308_),
    .B1(_05305_),
    .Y(_05340_));
 sky130_fd_sc_hd__a22o_1 _11555_ (.A1(_05218_),
    .A2(_05303_),
    .B1(_05339_),
    .B2(_05340_),
    .X(_05342_));
 sky130_fd_sc_hd__xnor2_1 _11556_ (.A(_05338_),
    .B(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__xnor2_1 _11557_ (.A(_05337_),
    .B(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__xnor2_1 _11558_ (.A(_05335_),
    .B(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__xnor2_1 _11559_ (.A(_05334_),
    .B(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__xnor2_1 _11560_ (.A(_05333_),
    .B(_05346_),
    .Y(_05347_));
 sky130_fd_sc_hd__o211a_1 _11561_ (.A1(_05329_),
    .A2(_05332_),
    .B1(_05347_),
    .C1(_05328_),
    .X(net124));
 sky130_fd_sc_hd__and2_1 _11562_ (.A(_02196_),
    .B(_03343_),
    .X(_05348_));
 sky130_fd_sc_hd__nor2_1 _11563_ (.A(_03354_),
    .B(_05348_),
    .Y(net128));
 sky130_fd_sc_hd__a22oi_1 _11564_ (.A1(net33),
    .A2(net12),
    .B1(net1),
    .B2(net44),
    .Y(_05349_));
 sky130_fd_sc_hd__nor2_1 _11565_ (.A(_00865_),
    .B(_05349_),
    .Y(net76));
 sky130_fd_sc_hd__nor2_1 _11566_ (.A(_00844_),
    .B(_00865_),
    .Y(_05351_));
 sky130_fd_sc_hd__nor2_1 _11567_ (.A(_00876_),
    .B(_05351_),
    .Y(net87));
 sky130_fd_sc_hd__nor2_1 _11568_ (.A(_00822_),
    .B(_00876_),
    .Y(_05352_));
 sky130_fd_sc_hd__nor2_1 _11569_ (.A(_00887_),
    .B(_05352_),
    .Y(net98));
 sky130_fd_sc_hd__a21o_1 _11570_ (.A1(_00789_),
    .A2(_00800_),
    .B1(_00887_),
    .X(_05353_));
 sky130_fd_sc_hd__and2_1 _11571_ (.A(_00898_),
    .B(_05353_),
    .X(net109));
 sky130_fd_sc_hd__buf_12 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_12 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_12 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_12 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_12 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_12 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_12 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_12 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_12 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_12 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_12 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_12 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_12 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_12 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_12 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_12 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_12 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_12 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_12 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_12 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_12 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_12 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_12 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_12 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_12 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_12 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_12 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_12 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_12 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_12 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_12 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_12 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_12 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_12 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_12 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_12 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_12 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_12 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_12 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_12 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_12 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_12 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_12 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_12 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_12 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_12 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_12 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_12 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_12 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_12 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_12 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_12 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_12 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_16 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_12 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_12 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_12 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_12 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_12 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_12 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_12 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_12 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_12 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_16 output65 (.A(net65),
    .X(result[0]));
 sky130_fd_sc_hd__clkbuf_16 output66 (.A(net66),
    .X(result[10]));
 sky130_fd_sc_hd__clkbuf_16 output67 (.A(net67),
    .X(result[11]));
 sky130_fd_sc_hd__clkbuf_16 output68 (.A(net68),
    .X(result[12]));
 sky130_fd_sc_hd__clkbuf_16 output69 (.A(net69),
    .X(result[13]));
 sky130_fd_sc_hd__clkbuf_16 output70 (.A(net70),
    .X(result[14]));
 sky130_fd_sc_hd__clkbuf_16 output71 (.A(net71),
    .X(result[15]));
 sky130_fd_sc_hd__clkbuf_16 output72 (.A(net72),
    .X(result[16]));
 sky130_fd_sc_hd__clkbuf_16 output73 (.A(net73),
    .X(result[17]));
 sky130_fd_sc_hd__clkbuf_16 output74 (.A(net74),
    .X(result[18]));
 sky130_fd_sc_hd__clkbuf_16 output75 (.A(net75),
    .X(result[19]));
 sky130_fd_sc_hd__clkbuf_16 output76 (.A(net76),
    .X(result[1]));
 sky130_fd_sc_hd__clkbuf_16 output77 (.A(net77),
    .X(result[20]));
 sky130_fd_sc_hd__clkbuf_16 output78 (.A(net78),
    .X(result[21]));
 sky130_fd_sc_hd__clkbuf_16 output79 (.A(net79),
    .X(result[22]));
 sky130_fd_sc_hd__clkbuf_16 output80 (.A(net80),
    .X(result[23]));
 sky130_fd_sc_hd__clkbuf_16 output81 (.A(net81),
    .X(result[24]));
 sky130_fd_sc_hd__clkbuf_16 output82 (.A(net82),
    .X(result[25]));
 sky130_fd_sc_hd__clkbuf_16 output83 (.A(net83),
    .X(result[26]));
 sky130_fd_sc_hd__clkbuf_16 output84 (.A(net84),
    .X(result[27]));
 sky130_fd_sc_hd__clkbuf_16 output85 (.A(net85),
    .X(result[28]));
 sky130_fd_sc_hd__clkbuf_16 output86 (.A(net86),
    .X(result[29]));
 sky130_fd_sc_hd__clkbuf_16 output87 (.A(net87),
    .X(result[2]));
 sky130_fd_sc_hd__clkbuf_16 output88 (.A(net88),
    .X(result[30]));
 sky130_fd_sc_hd__clkbuf_16 output89 (.A(net89),
    .X(result[31]));
 sky130_fd_sc_hd__clkbuf_16 output90 (.A(net90),
    .X(result[32]));
 sky130_fd_sc_hd__clkbuf_16 output91 (.A(net91),
    .X(result[33]));
 sky130_fd_sc_hd__clkbuf_16 output92 (.A(net92),
    .X(result[34]));
 sky130_fd_sc_hd__clkbuf_16 output93 (.A(net93),
    .X(result[35]));
 sky130_fd_sc_hd__clkbuf_16 output94 (.A(net94),
    .X(result[36]));
 sky130_fd_sc_hd__clkbuf_16 output95 (.A(net95),
    .X(result[37]));
 sky130_fd_sc_hd__clkbuf_16 output96 (.A(net96),
    .X(result[38]));
 sky130_fd_sc_hd__clkbuf_16 output97 (.A(net97),
    .X(result[39]));
 sky130_fd_sc_hd__clkbuf_16 output98 (.A(net98),
    .X(result[3]));
 sky130_fd_sc_hd__clkbuf_16 output99 (.A(net99),
    .X(result[40]));
 sky130_fd_sc_hd__clkbuf_16 output100 (.A(net100),
    .X(result[41]));
 sky130_fd_sc_hd__clkbuf_16 output101 (.A(net101),
    .X(result[42]));
 sky130_fd_sc_hd__clkbuf_16 output102 (.A(net102),
    .X(result[43]));
 sky130_fd_sc_hd__clkbuf_16 output103 (.A(net103),
    .X(result[44]));
 sky130_fd_sc_hd__clkbuf_16 output104 (.A(net104),
    .X(result[45]));
 sky130_fd_sc_hd__clkbuf_16 output105 (.A(net105),
    .X(result[46]));
 sky130_fd_sc_hd__clkbuf_16 output106 (.A(net106),
    .X(result[47]));
 sky130_fd_sc_hd__clkbuf_16 output107 (.A(net107),
    .X(result[48]));
 sky130_fd_sc_hd__clkbuf_16 output108 (.A(net108),
    .X(result[49]));
 sky130_fd_sc_hd__clkbuf_16 output109 (.A(net109),
    .X(result[4]));
 sky130_fd_sc_hd__clkbuf_16 output110 (.A(net110),
    .X(result[50]));
 sky130_fd_sc_hd__clkbuf_16 output111 (.A(net111),
    .X(result[51]));
 sky130_fd_sc_hd__clkbuf_16 output112 (.A(net112),
    .X(result[52]));
 sky130_fd_sc_hd__clkbuf_16 output113 (.A(net113),
    .X(result[53]));
 sky130_fd_sc_hd__clkbuf_16 output114 (.A(net114),
    .X(result[54]));
 sky130_fd_sc_hd__clkbuf_16 output115 (.A(net115),
    .X(result[55]));
 sky130_fd_sc_hd__clkbuf_16 output116 (.A(net116),
    .X(result[56]));
 sky130_fd_sc_hd__clkbuf_16 output117 (.A(net117),
    .X(result[57]));
 sky130_fd_sc_hd__clkbuf_16 output118 (.A(net118),
    .X(result[58]));
 sky130_fd_sc_hd__clkbuf_16 output119 (.A(net119),
    .X(result[59]));
 sky130_fd_sc_hd__clkbuf_16 output120 (.A(net120),
    .X(result[5]));
 sky130_fd_sc_hd__clkbuf_16 output121 (.A(net121),
    .X(result[60]));
 sky130_fd_sc_hd__clkbuf_16 output122 (.A(net122),
    .X(result[61]));
 sky130_fd_sc_hd__clkbuf_16 output123 (.A(net123),
    .X(result[62]));
 sky130_fd_sc_hd__clkbuf_16 output124 (.A(net124),
    .X(result[63]));
 sky130_fd_sc_hd__clkbuf_16 output125 (.A(net125),
    .X(result[6]));
 sky130_fd_sc_hd__clkbuf_16 output126 (.A(net126),
    .X(result[7]));
 sky130_fd_sc_hd__clkbuf_16 output127 (.A(net127),
    .X(result[8]));
 sky130_fd_sc_hd__clkbuf_16 output128 (.A(net128),
    .X(result[9]));
endmodule
