module tree_multiplier_route (A,
    B,
    z);
 input [31:0] A;
 input [31:0] B;
 output [63:0] z;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire \genblk2[10].rca.ripple_adders[0].fa.a ;
 wire \genblk2[10].rca.ripple_adders[10].fa.a ;
 wire \genblk2[10].rca.ripple_adders[11].fa.sum ;
 wire \genblk2[10].rca.ripple_adders[1].fa.a ;
 wire \genblk2[10].rca.ripple_adders[2].fa.a ;
 wire \genblk2[10].rca.ripple_adders[3].fa.a ;
 wire \genblk2[10].rca.ripple_adders[4].fa.a ;
 wire \genblk2[10].rca.ripple_adders[5].fa.a ;
 wire \genblk2[10].rca.ripple_adders[6].fa.a ;
 wire \genblk2[10].rca.ripple_adders[7].fa.a ;
 wire \genblk2[10].rca.ripple_adders[8].fa.a ;
 wire \genblk2[10].rca.ripple_adders[9].fa.a ;
 wire \genblk2[11].rca.ripple_adders[12].fa.sum ;
 wire \genblk2[12].rca.ripple_adders[13].fa.sum ;
 wire \genblk2[13].rca.ripple_adders[14].fa.sum ;
 wire \genblk2[14].rca.ripple_adders[15].fa.sum ;
 wire \genblk2[15].rca.ripple_adders[16].fa.sum ;
 wire \genblk2[16].rca.ripple_adders[17].fa.sum ;
 wire \genblk2[17].rca.ripple_adders[18].fa.sum ;
 wire \genblk2[18].rca.ripple_adders[19].fa.sum ;
 wire \genblk2[19].rca.ripple_adders[20].fa.sum ;
 wire \genblk2[20].rca.ripple_adders[21].fa.sum ;
 wire \genblk2[21].rca.ripple_adders[22].fa.sum ;
 wire \genblk2[22].rca.ripple_adders[23].fa.sum ;
 wire \genblk2[23].rca.ripple_adders[24].fa.sum ;
 wire \genblk2[24].rca.ripple_adders[25].fa.sum ;
 wire \genblk2[25].rca.ripple_adders[26].fa.sum ;
 wire \genblk2[26].rca.ripple_adders[27].fa.sum ;
 wire \genblk2[27].rca.ripple_adders[28].fa.sum ;
 wire \genblk2[28].rca.ripple_adders[29].fa.sum ;
 wire \genblk2[29].rca.ripple_adders[30].fa.sum ;
 wire \genblk2[30].rca.ripple_adders[31].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[0].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[10].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[11].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[12].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[13].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[14].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[15].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[16].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[17].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[18].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[19].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[1].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[20].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[21].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[22].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[23].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[24].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[25].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[26].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[27].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[28].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[29].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[2].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[30].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[31].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[3].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[4].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[5].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[6].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[7].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[8].fa.sum ;
 wire \genblk2[30].rca1.ripple_adders[9].fa.sum ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;

 sky130_fd_sc_hd__nand2_1 _04984_ (.A(net1),
    .B(net55),
    .Y(_00287_));
 sky130_fd_sc_hd__nand2_1 _04985_ (.A(net23),
    .B(net33),
    .Y(_00298_));
 sky130_fd_sc_hd__nand2_1 _04986_ (.A(net1),
    .B(net33),
    .Y(_00309_));
 sky130_fd_sc_hd__inv_2 _04987_ (.A(_00309_),
    .Y(\genblk2[10].rca.ripple_adders[0].fa.a ));
 sky130_fd_sc_hd__a31o_1 _04988_ (.A1(net12),
    .A2(net44),
    .A3(_00309_),
    .B1(_00298_),
    .X(_00329_));
 sky130_fd_sc_hd__nand4_1 _04989_ (.A(net12),
    .B(net44),
    .C(_00298_),
    .D(_00309_),
    .Y(_00340_));
 sky130_fd_sc_hd__a21oi_1 _04990_ (.A1(_00329_),
    .A2(_00340_),
    .B1(_00287_),
    .Y(_00351_));
 sky130_fd_sc_hd__a22o_1 _04991_ (.A1(net26),
    .A2(net33),
    .B1(net44),
    .B2(net23),
    .X(_00362_));
 sky130_fd_sc_hd__nand4_1 _04992_ (.A(net26),
    .B(net23),
    .C(net33),
    .D(net44),
    .Y(_00373_));
 sky130_fd_sc_hd__nand2_4 _04993_ (.A(net33),
    .B(net44),
    .Y(_00384_));
 sky130_fd_sc_hd__nand2_1 _04994_ (.A(net12),
    .B(net1),
    .Y(_00395_));
 sky130_fd_sc_hd__o2111a_1 _04995_ (.A1(net23),
    .A2(net1),
    .B1(net33),
    .C1(net44),
    .D1(net12),
    .X(_00406_));
 sky130_fd_sc_hd__nand3_1 _04996_ (.A(_00362_),
    .B(_00373_),
    .C(_00406_),
    .Y(_00417_));
 sky130_fd_sc_hd__a21o_1 _04997_ (.A1(_00362_),
    .A2(_00373_),
    .B1(_00406_),
    .X(_00428_));
 sky130_fd_sc_hd__and4_1 _04998_ (.A(net12),
    .B(net55),
    .C(_00417_),
    .D(_00428_),
    .X(_00439_));
 sky130_fd_sc_hd__a22o_1 _04999_ (.A1(net12),
    .A2(net55),
    .B1(_00417_),
    .B2(_00428_),
    .X(_00450_));
 sky130_fd_sc_hd__nand2b_1 _05000_ (.A_N(_00439_),
    .B(_00450_),
    .Y(_00460_));
 sky130_fd_sc_hd__xnor2_1 _05001_ (.A(_00351_),
    .B(_00460_),
    .Y(_00471_));
 sky130_fd_sc_hd__and3_1 _05002_ (.A(net1),
    .B(net58),
    .C(_00471_),
    .X(_00482_));
 sky130_fd_sc_hd__a21o_1 _05003_ (.A1(_00351_),
    .A2(_00450_),
    .B1(_00439_),
    .X(_00493_));
 sky130_fd_sc_hd__a21bo_1 _05004_ (.A1(_00362_),
    .A2(_00406_),
    .B1_N(_00373_),
    .X(_00504_));
 sky130_fd_sc_hd__and4_1 _05005_ (.A(net26),
    .B(net33),
    .C(net44),
    .D(net27),
    .X(_00515_));
 sky130_fd_sc_hd__a22o_1 _05006_ (.A1(net26),
    .A2(net44),
    .B1(net27),
    .B2(net33),
    .X(_00526_));
 sky130_fd_sc_hd__nand2b_1 _05007_ (.A_N(_00515_),
    .B(_00526_),
    .Y(_00537_));
 sky130_fd_sc_hd__xnor2_1 _05008_ (.A(_00504_),
    .B(_00537_),
    .Y(_00548_));
 sky130_fd_sc_hd__nand2_1 _05009_ (.A(net23),
    .B(net55),
    .Y(_00559_));
 sky130_fd_sc_hd__and3_1 _05010_ (.A(net23),
    .B(net55),
    .C(_00548_),
    .X(_00570_));
 sky130_fd_sc_hd__xnor2_1 _05011_ (.A(_00548_),
    .B(_00559_),
    .Y(_00580_));
 sky130_fd_sc_hd__xor2_1 _05012_ (.A(_00493_),
    .B(_00580_),
    .X(_00591_));
 sky130_fd_sc_hd__and3_1 _05013_ (.A(net12),
    .B(net58),
    .C(_00591_),
    .X(_00602_));
 sky130_fd_sc_hd__a21o_1 _05014_ (.A1(net12),
    .A2(net58),
    .B1(_00591_),
    .X(_00613_));
 sky130_fd_sc_hd__nand2b_1 _05015_ (.A_N(_00602_),
    .B(_00613_),
    .Y(_00624_));
 sky130_fd_sc_hd__xnor2_1 _05016_ (.A(_00482_),
    .B(_00624_),
    .Y(_00635_));
 sky130_fd_sc_hd__and3_1 _05017_ (.A(net1),
    .B(net59),
    .C(_00635_),
    .X(_00646_));
 sky130_fd_sc_hd__a21o_1 _05018_ (.A1(_00482_),
    .A2(_00613_),
    .B1(_00602_),
    .X(_00657_));
 sky130_fd_sc_hd__a21o_1 _05019_ (.A1(_00493_),
    .A2(_00580_),
    .B1(_00570_),
    .X(_00668_));
 sky130_fd_sc_hd__and4_1 _05020_ (.A(net33),
    .B(net44),
    .C(net28),
    .D(net27),
    .X(_00679_));
 sky130_fd_sc_hd__a22o_1 _05021_ (.A1(net33),
    .A2(net28),
    .B1(net27),
    .B2(net44),
    .X(_00690_));
 sky130_fd_sc_hd__nand2b_1 _05022_ (.A_N(_00679_),
    .B(_00690_),
    .Y(_00701_));
 sky130_fd_sc_hd__a21o_1 _05023_ (.A1(_00504_),
    .A2(_00526_),
    .B1(_00515_),
    .X(_00712_));
 sky130_fd_sc_hd__xnor2_1 _05024_ (.A(_00701_),
    .B(_00712_),
    .Y(_00722_));
 sky130_fd_sc_hd__nand2_1 _05025_ (.A(net26),
    .B(net55),
    .Y(_00733_));
 sky130_fd_sc_hd__and3_1 _05026_ (.A(net26),
    .B(net55),
    .C(_00722_),
    .X(_00744_));
 sky130_fd_sc_hd__nand2b_1 _05027_ (.A_N(_00722_),
    .B(_00733_),
    .Y(_00755_));
 sky130_fd_sc_hd__xor2_1 _05028_ (.A(_00722_),
    .B(_00733_),
    .X(_00766_));
 sky130_fd_sc_hd__xnor2_1 _05029_ (.A(_00668_),
    .B(_00766_),
    .Y(_00777_));
 sky130_fd_sc_hd__nand2_1 _05030_ (.A(net23),
    .B(net58),
    .Y(_00788_));
 sky130_fd_sc_hd__and3_1 _05031_ (.A(net23),
    .B(net58),
    .C(_00777_),
    .X(_00799_));
 sky130_fd_sc_hd__xnor2_1 _05032_ (.A(_00777_),
    .B(_00788_),
    .Y(_00810_));
 sky130_fd_sc_hd__xor2_1 _05033_ (.A(_00657_),
    .B(_00810_),
    .X(_00821_));
 sky130_fd_sc_hd__and3_1 _05034_ (.A(net12),
    .B(net59),
    .C(_00821_),
    .X(_00832_));
 sky130_fd_sc_hd__a21o_1 _05035_ (.A1(net12),
    .A2(net59),
    .B1(_00821_),
    .X(_00843_));
 sky130_fd_sc_hd__nand2b_1 _05036_ (.A_N(_00832_),
    .B(_00843_),
    .Y(_00853_));
 sky130_fd_sc_hd__xnor2_1 _05037_ (.A(_00646_),
    .B(_00853_),
    .Y(_00864_));
 sky130_fd_sc_hd__and3_1 _05038_ (.A(net1),
    .B(net60),
    .C(_00864_),
    .X(_00875_));
 sky130_fd_sc_hd__a21o_1 _05039_ (.A1(_00646_),
    .A2(_00843_),
    .B1(_00832_),
    .X(_00886_));
 sky130_fd_sc_hd__a21o_1 _05040_ (.A1(_00657_),
    .A2(_00810_),
    .B1(_00799_),
    .X(_00897_));
 sky130_fd_sc_hd__a21o_1 _05041_ (.A1(_00668_),
    .A2(_00755_),
    .B1(_00744_),
    .X(_00908_));
 sky130_fd_sc_hd__and4_1 _05042_ (.A(net33),
    .B(net44),
    .C(net29),
    .D(net28),
    .X(_00919_));
 sky130_fd_sc_hd__a22o_1 _05043_ (.A1(net33),
    .A2(net29),
    .B1(net28),
    .B2(net44),
    .X(_00930_));
 sky130_fd_sc_hd__nand2b_1 _05044_ (.A_N(_00919_),
    .B(_00930_),
    .Y(_00941_));
 sky130_fd_sc_hd__a21o_1 _05045_ (.A1(_00690_),
    .A2(_00712_),
    .B1(_00679_),
    .X(_00952_));
 sky130_fd_sc_hd__xnor2_1 _05046_ (.A(_00941_),
    .B(_00952_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2_1 _05047_ (.A(net55),
    .B(net27),
    .Y(_00974_));
 sky130_fd_sc_hd__and3_1 _05048_ (.A(net55),
    .B(net27),
    .C(_00963_),
    .X(_00985_));
 sky130_fd_sc_hd__nand2b_1 _05049_ (.A_N(_00963_),
    .B(_00974_),
    .Y(_00996_));
 sky130_fd_sc_hd__xor2_1 _05050_ (.A(_00963_),
    .B(_00974_),
    .X(_01006_));
 sky130_fd_sc_hd__xnor2_1 _05051_ (.A(_00908_),
    .B(_01006_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _05052_ (.A(net26),
    .B(net58),
    .Y(_01028_));
 sky130_fd_sc_hd__and3_1 _05053_ (.A(net26),
    .B(net58),
    .C(_01017_),
    .X(_01039_));
 sky130_fd_sc_hd__xnor2_1 _05054_ (.A(_01017_),
    .B(_01028_),
    .Y(_01050_));
 sky130_fd_sc_hd__xor2_1 _05055_ (.A(_00897_),
    .B(_01050_),
    .X(_01061_));
 sky130_fd_sc_hd__nand2_1 _05056_ (.A(net23),
    .B(net59),
    .Y(_01072_));
 sky130_fd_sc_hd__and3_1 _05057_ (.A(net23),
    .B(net59),
    .C(_01061_),
    .X(_01083_));
 sky130_fd_sc_hd__xnor2_1 _05058_ (.A(_01061_),
    .B(_01072_),
    .Y(_01094_));
 sky130_fd_sc_hd__xor2_1 _05059_ (.A(_00886_),
    .B(_01094_),
    .X(_01105_));
 sky130_fd_sc_hd__and3_1 _05060_ (.A(net12),
    .B(net60),
    .C(_01105_),
    .X(_01116_));
 sky130_fd_sc_hd__a21o_1 _05061_ (.A1(net12),
    .A2(net60),
    .B1(_01105_),
    .X(_01127_));
 sky130_fd_sc_hd__nand2b_1 _05062_ (.A_N(_01116_),
    .B(_01127_),
    .Y(_01138_));
 sky130_fd_sc_hd__xnor2_1 _05063_ (.A(_00875_),
    .B(_01138_),
    .Y(_01149_));
 sky130_fd_sc_hd__and3_1 _05064_ (.A(net1),
    .B(net61),
    .C(_01149_),
    .X(_01159_));
 sky130_fd_sc_hd__a21o_1 _05065_ (.A1(_00875_),
    .A2(_01127_),
    .B1(_01116_),
    .X(_01170_));
 sky130_fd_sc_hd__a21o_1 _05066_ (.A1(_00886_),
    .A2(_01094_),
    .B1(_01083_),
    .X(_01181_));
 sky130_fd_sc_hd__a21o_1 _05067_ (.A1(_00897_),
    .A2(_01050_),
    .B1(_01039_),
    .X(_01192_));
 sky130_fd_sc_hd__a21o_1 _05068_ (.A1(_00908_),
    .A2(_00996_),
    .B1(_00985_),
    .X(_01203_));
 sky130_fd_sc_hd__and4_1 _05069_ (.A(net33),
    .B(net44),
    .C(net30),
    .D(net29),
    .X(_01214_));
 sky130_fd_sc_hd__a22o_1 _05070_ (.A1(net33),
    .A2(net30),
    .B1(net29),
    .B2(net44),
    .X(_01225_));
 sky130_fd_sc_hd__nand2b_1 _05071_ (.A_N(_01214_),
    .B(_01225_),
    .Y(_01236_));
 sky130_fd_sc_hd__a21o_1 _05072_ (.A1(_00930_),
    .A2(_00952_),
    .B1(_00919_),
    .X(_01247_));
 sky130_fd_sc_hd__xnor2_1 _05073_ (.A(_01236_),
    .B(_01247_),
    .Y(_01258_));
 sky130_fd_sc_hd__nand2_1 _05074_ (.A(net55),
    .B(net28),
    .Y(_01269_));
 sky130_fd_sc_hd__and3_1 _05075_ (.A(net55),
    .B(net28),
    .C(_01258_),
    .X(_01280_));
 sky130_fd_sc_hd__nand2b_1 _05076_ (.A_N(_01258_),
    .B(_01269_),
    .Y(_01291_));
 sky130_fd_sc_hd__xor2_1 _05077_ (.A(_01258_),
    .B(_01269_),
    .X(_01302_));
 sky130_fd_sc_hd__xnor2_1 _05078_ (.A(_01203_),
    .B(_01302_),
    .Y(_01312_));
 sky130_fd_sc_hd__nand2_1 _05079_ (.A(net58),
    .B(net27),
    .Y(_01323_));
 sky130_fd_sc_hd__and3_1 _05080_ (.A(net58),
    .B(net27),
    .C(_01312_),
    .X(_01334_));
 sky130_fd_sc_hd__xnor2_1 _05081_ (.A(_01312_),
    .B(_01323_),
    .Y(_01345_));
 sky130_fd_sc_hd__xor2_1 _05082_ (.A(_01192_),
    .B(_01345_),
    .X(_01356_));
 sky130_fd_sc_hd__nand2_1 _05083_ (.A(net26),
    .B(net59),
    .Y(_01367_));
 sky130_fd_sc_hd__and3_1 _05084_ (.A(net26),
    .B(net59),
    .C(_01356_),
    .X(_01378_));
 sky130_fd_sc_hd__xnor2_1 _05085_ (.A(_01356_),
    .B(_01367_),
    .Y(_01389_));
 sky130_fd_sc_hd__xor2_1 _05086_ (.A(_01181_),
    .B(_01389_),
    .X(_01400_));
 sky130_fd_sc_hd__nand2_1 _05087_ (.A(net23),
    .B(net60),
    .Y(_01411_));
 sky130_fd_sc_hd__and3_1 _05088_ (.A(net23),
    .B(net60),
    .C(_01400_),
    .X(_01422_));
 sky130_fd_sc_hd__xnor2_1 _05089_ (.A(_01400_),
    .B(_01411_),
    .Y(_01433_));
 sky130_fd_sc_hd__xor2_1 _05090_ (.A(_01170_),
    .B(_01433_),
    .X(_01444_));
 sky130_fd_sc_hd__and3_1 _05091_ (.A(net12),
    .B(net61),
    .C(_01444_),
    .X(_01455_));
 sky130_fd_sc_hd__a21o_1 _05092_ (.A1(net12),
    .A2(net61),
    .B1(_01444_),
    .X(_01466_));
 sky130_fd_sc_hd__nand2b_1 _05093_ (.A_N(_01455_),
    .B(_01466_),
    .Y(_01476_));
 sky130_fd_sc_hd__xnor2_1 _05094_ (.A(_01159_),
    .B(_01476_),
    .Y(_01487_));
 sky130_fd_sc_hd__and3_1 _05095_ (.A(net1),
    .B(net62),
    .C(_01487_),
    .X(_01498_));
 sky130_fd_sc_hd__a21o_1 _05096_ (.A1(_01159_),
    .A2(_01466_),
    .B1(_01455_),
    .X(_01509_));
 sky130_fd_sc_hd__a21o_1 _05097_ (.A1(_01170_),
    .A2(_01433_),
    .B1(_01422_),
    .X(_01520_));
 sky130_fd_sc_hd__a21o_1 _05098_ (.A1(_01181_),
    .A2(_01389_),
    .B1(_01378_),
    .X(_01531_));
 sky130_fd_sc_hd__a21o_1 _05099_ (.A1(_01192_),
    .A2(_01345_),
    .B1(_01334_),
    .X(_01542_));
 sky130_fd_sc_hd__a21o_1 _05100_ (.A1(_01203_),
    .A2(_01291_),
    .B1(_01280_),
    .X(_01553_));
 sky130_fd_sc_hd__and4_1 _05101_ (.A(net33),
    .B(net44),
    .C(net31),
    .D(net30),
    .X(_01564_));
 sky130_fd_sc_hd__a22o_1 _05102_ (.A1(net33),
    .A2(net31),
    .B1(net30),
    .B2(net44),
    .X(_01575_));
 sky130_fd_sc_hd__nand2b_1 _05103_ (.A_N(_01564_),
    .B(_01575_),
    .Y(_01586_));
 sky130_fd_sc_hd__a21o_1 _05104_ (.A1(_01225_),
    .A2(_01247_),
    .B1(_01214_),
    .X(_01597_));
 sky130_fd_sc_hd__xnor2_1 _05105_ (.A(_01586_),
    .B(_01597_),
    .Y(_01608_));
 sky130_fd_sc_hd__nand2_1 _05106_ (.A(net55),
    .B(net29),
    .Y(_01619_));
 sky130_fd_sc_hd__and3_1 _05107_ (.A(net55),
    .B(net29),
    .C(_01608_),
    .X(_01630_));
 sky130_fd_sc_hd__nand2b_1 _05108_ (.A_N(_01608_),
    .B(_01619_),
    .Y(_01640_));
 sky130_fd_sc_hd__xor2_1 _05109_ (.A(_01608_),
    .B(_01619_),
    .X(_01651_));
 sky130_fd_sc_hd__xnor2_1 _05110_ (.A(_01553_),
    .B(_01651_),
    .Y(_01662_));
 sky130_fd_sc_hd__nand2_1 _05111_ (.A(net58),
    .B(net28),
    .Y(_01673_));
 sky130_fd_sc_hd__and3_1 _05112_ (.A(net58),
    .B(net28),
    .C(_01662_),
    .X(_01684_));
 sky130_fd_sc_hd__xnor2_1 _05113_ (.A(_01662_),
    .B(_01673_),
    .Y(_01695_));
 sky130_fd_sc_hd__xor2_1 _05114_ (.A(_01542_),
    .B(_01695_),
    .X(_01706_));
 sky130_fd_sc_hd__nand2_1 _05115_ (.A(net59),
    .B(net27),
    .Y(_01717_));
 sky130_fd_sc_hd__and3_1 _05116_ (.A(net59),
    .B(net27),
    .C(_01706_),
    .X(_01728_));
 sky130_fd_sc_hd__xnor2_1 _05117_ (.A(_01706_),
    .B(_01717_),
    .Y(_01739_));
 sky130_fd_sc_hd__xor2_1 _05118_ (.A(_01531_),
    .B(_01739_),
    .X(_01750_));
 sky130_fd_sc_hd__nand2_1 _05119_ (.A(net26),
    .B(net60),
    .Y(_01761_));
 sky130_fd_sc_hd__and3_1 _05120_ (.A(net26),
    .B(net60),
    .C(_01750_),
    .X(_01772_));
 sky130_fd_sc_hd__xnor2_1 _05121_ (.A(_01750_),
    .B(_01761_),
    .Y(_01783_));
 sky130_fd_sc_hd__xor2_1 _05122_ (.A(_01520_),
    .B(_01783_),
    .X(_01794_));
 sky130_fd_sc_hd__nand2_1 _05123_ (.A(net23),
    .B(net61),
    .Y(_01805_));
 sky130_fd_sc_hd__and3_1 _05124_ (.A(net23),
    .B(net61),
    .C(_01794_),
    .X(_01816_));
 sky130_fd_sc_hd__xnor2_1 _05125_ (.A(_01794_),
    .B(_01805_),
    .Y(_01827_));
 sky130_fd_sc_hd__xor2_1 _05126_ (.A(_01509_),
    .B(_01827_),
    .X(_01838_));
 sky130_fd_sc_hd__and3_1 _05127_ (.A(net12),
    .B(net62),
    .C(_01838_),
    .X(_01849_));
 sky130_fd_sc_hd__a21o_1 _05128_ (.A1(net12),
    .A2(net62),
    .B1(_01838_),
    .X(_01860_));
 sky130_fd_sc_hd__nand2b_1 _05129_ (.A_N(_01849_),
    .B(_01860_),
    .Y(_01871_));
 sky130_fd_sc_hd__xnor2_1 _05130_ (.A(_01498_),
    .B(_01871_),
    .Y(_01882_));
 sky130_fd_sc_hd__and3_1 _05131_ (.A(net1),
    .B(net63),
    .C(_01882_),
    .X(_01893_));
 sky130_fd_sc_hd__a21o_1 _05132_ (.A1(_01498_),
    .A2(_01860_),
    .B1(_01849_),
    .X(_01904_));
 sky130_fd_sc_hd__a21o_1 _05133_ (.A1(_01509_),
    .A2(_01827_),
    .B1(_01816_),
    .X(_01915_));
 sky130_fd_sc_hd__a21o_1 _05134_ (.A1(_01520_),
    .A2(_01783_),
    .B1(_01772_),
    .X(_01926_));
 sky130_fd_sc_hd__a21o_1 _05135_ (.A1(_01531_),
    .A2(_01739_),
    .B1(_01728_),
    .X(_01937_));
 sky130_fd_sc_hd__a21o_1 _05136_ (.A1(_01542_),
    .A2(_01695_),
    .B1(_01684_),
    .X(_01948_));
 sky130_fd_sc_hd__a21o_1 _05137_ (.A1(_01553_),
    .A2(_01640_),
    .B1(_01630_),
    .X(_01959_));
 sky130_fd_sc_hd__and4_1 _05138_ (.A(net33),
    .B(net44),
    .C(net32),
    .D(net31),
    .X(_01970_));
 sky130_fd_sc_hd__a22o_1 _05139_ (.A1(net33),
    .A2(net32),
    .B1(net31),
    .B2(net44),
    .X(_01981_));
 sky130_fd_sc_hd__nand2b_1 _05140_ (.A_N(_01970_),
    .B(_01981_),
    .Y(_01992_));
 sky130_fd_sc_hd__a21o_1 _05141_ (.A1(_01575_),
    .A2(_01597_),
    .B1(_01564_),
    .X(_02003_));
 sky130_fd_sc_hd__xnor2_1 _05142_ (.A(_01992_),
    .B(_02003_),
    .Y(_02014_));
 sky130_fd_sc_hd__nand2_1 _05143_ (.A(net55),
    .B(net30),
    .Y(_02025_));
 sky130_fd_sc_hd__and3_1 _05144_ (.A(net55),
    .B(net30),
    .C(_02014_),
    .X(_02036_));
 sky130_fd_sc_hd__nand2b_1 _05145_ (.A_N(_02014_),
    .B(_02025_),
    .Y(_02047_));
 sky130_fd_sc_hd__xor2_1 _05146_ (.A(_02014_),
    .B(_02025_),
    .X(_02058_));
 sky130_fd_sc_hd__xnor2_1 _05147_ (.A(_01959_),
    .B(_02058_),
    .Y(_02069_));
 sky130_fd_sc_hd__nand2_1 _05148_ (.A(net58),
    .B(net29),
    .Y(_02080_));
 sky130_fd_sc_hd__and3_1 _05149_ (.A(net58),
    .B(net29),
    .C(_02069_),
    .X(_02091_));
 sky130_fd_sc_hd__xnor2_1 _05150_ (.A(_02069_),
    .B(_02080_),
    .Y(_02102_));
 sky130_fd_sc_hd__xor2_1 _05151_ (.A(_01948_),
    .B(_02102_),
    .X(_02113_));
 sky130_fd_sc_hd__nand2_1 _05152_ (.A(net59),
    .B(net28),
    .Y(_02124_));
 sky130_fd_sc_hd__and3_1 _05153_ (.A(net59),
    .B(net28),
    .C(_02113_),
    .X(_02135_));
 sky130_fd_sc_hd__xnor2_1 _05154_ (.A(_02113_),
    .B(_02124_),
    .Y(_02146_));
 sky130_fd_sc_hd__xor2_1 _05155_ (.A(_01937_),
    .B(_02146_),
    .X(_02157_));
 sky130_fd_sc_hd__nand2_1 _05156_ (.A(net60),
    .B(net27),
    .Y(_02168_));
 sky130_fd_sc_hd__and3_1 _05157_ (.A(net60),
    .B(net27),
    .C(_02157_),
    .X(_02179_));
 sky130_fd_sc_hd__xnor2_1 _05158_ (.A(_02157_),
    .B(_02168_),
    .Y(_02190_));
 sky130_fd_sc_hd__xor2_1 _05159_ (.A(_01926_),
    .B(_02190_),
    .X(_02201_));
 sky130_fd_sc_hd__nand2_1 _05160_ (.A(net26),
    .B(net61),
    .Y(_02212_));
 sky130_fd_sc_hd__and3_1 _05161_ (.A(net26),
    .B(net61),
    .C(_02201_),
    .X(_02223_));
 sky130_fd_sc_hd__xnor2_1 _05162_ (.A(_02201_),
    .B(_02212_),
    .Y(_02234_));
 sky130_fd_sc_hd__xor2_1 _05163_ (.A(_01915_),
    .B(_02234_),
    .X(_02245_));
 sky130_fd_sc_hd__nand2_1 _05164_ (.A(net23),
    .B(net62),
    .Y(_02256_));
 sky130_fd_sc_hd__and3_1 _05165_ (.A(net23),
    .B(net62),
    .C(_02245_),
    .X(_02267_));
 sky130_fd_sc_hd__xnor2_1 _05166_ (.A(_02245_),
    .B(_02256_),
    .Y(_02278_));
 sky130_fd_sc_hd__xor2_1 _05167_ (.A(_01904_),
    .B(_02278_),
    .X(_02289_));
 sky130_fd_sc_hd__and3_1 _05168_ (.A(net12),
    .B(net63),
    .C(_02289_),
    .X(_02300_));
 sky130_fd_sc_hd__a21o_1 _05169_ (.A1(net12),
    .A2(net63),
    .B1(_02289_),
    .X(_02311_));
 sky130_fd_sc_hd__nand2b_1 _05170_ (.A_N(_02300_),
    .B(_02311_),
    .Y(_02322_));
 sky130_fd_sc_hd__xnor2_1 _05171_ (.A(_01893_),
    .B(_02322_),
    .Y(_02333_));
 sky130_fd_sc_hd__and3_1 _05172_ (.A(net64),
    .B(net1),
    .C(_02333_),
    .X(_02344_));
 sky130_fd_sc_hd__a21o_1 _05173_ (.A1(_01893_),
    .A2(_02311_),
    .B1(_02300_),
    .X(_02355_));
 sky130_fd_sc_hd__a21o_1 _05174_ (.A1(_01904_),
    .A2(_02278_),
    .B1(_02267_),
    .X(_02366_));
 sky130_fd_sc_hd__a21o_1 _05175_ (.A1(_01915_),
    .A2(_02234_),
    .B1(_02223_),
    .X(_02377_));
 sky130_fd_sc_hd__a21o_1 _05176_ (.A1(_01926_),
    .A2(_02190_),
    .B1(_02179_),
    .X(_02388_));
 sky130_fd_sc_hd__a21o_1 _05177_ (.A1(_01937_),
    .A2(_02146_),
    .B1(_02135_),
    .X(_02399_));
 sky130_fd_sc_hd__a21o_1 _05178_ (.A1(_01948_),
    .A2(_02102_),
    .B1(_02091_),
    .X(_02410_));
 sky130_fd_sc_hd__a21o_1 _05179_ (.A1(_01959_),
    .A2(_02047_),
    .B1(_02036_),
    .X(_02421_));
 sky130_fd_sc_hd__and4_1 _05180_ (.A(net33),
    .B(net44),
    .C(net2),
    .D(net32),
    .X(_02432_));
 sky130_fd_sc_hd__a22o_1 _05181_ (.A1(net33),
    .A2(net2),
    .B1(net32),
    .B2(net44),
    .X(_02443_));
 sky130_fd_sc_hd__nand2b_1 _05182_ (.A_N(_02432_),
    .B(_02443_),
    .Y(_02454_));
 sky130_fd_sc_hd__a21o_1 _05183_ (.A1(_01981_),
    .A2(_02003_),
    .B1(_01970_),
    .X(_02465_));
 sky130_fd_sc_hd__xnor2_1 _05184_ (.A(_02454_),
    .B(_02465_),
    .Y(_02476_));
 sky130_fd_sc_hd__nand2_1 _05185_ (.A(net55),
    .B(net31),
    .Y(_02487_));
 sky130_fd_sc_hd__and3_1 _05186_ (.A(net55),
    .B(net31),
    .C(_02476_),
    .X(_02498_));
 sky130_fd_sc_hd__nand2b_1 _05187_ (.A_N(_02476_),
    .B(_02487_),
    .Y(_02509_));
 sky130_fd_sc_hd__xor2_1 _05188_ (.A(_02476_),
    .B(_02487_),
    .X(_02520_));
 sky130_fd_sc_hd__xnor2_1 _05189_ (.A(_02421_),
    .B(_02520_),
    .Y(_02531_));
 sky130_fd_sc_hd__nand2_1 _05190_ (.A(net58),
    .B(net30),
    .Y(_02542_));
 sky130_fd_sc_hd__and3_1 _05191_ (.A(net58),
    .B(net30),
    .C(_02531_),
    .X(_02553_));
 sky130_fd_sc_hd__xnor2_1 _05192_ (.A(_02531_),
    .B(_02542_),
    .Y(_02564_));
 sky130_fd_sc_hd__xor2_1 _05193_ (.A(_02410_),
    .B(_02564_),
    .X(_02575_));
 sky130_fd_sc_hd__nand2_1 _05194_ (.A(net59),
    .B(net29),
    .Y(_02586_));
 sky130_fd_sc_hd__and3_1 _05195_ (.A(net59),
    .B(net29),
    .C(_02575_),
    .X(_02597_));
 sky130_fd_sc_hd__xnor2_1 _05196_ (.A(_02575_),
    .B(_02586_),
    .Y(_02608_));
 sky130_fd_sc_hd__xor2_1 _05197_ (.A(_02399_),
    .B(_02608_),
    .X(_02619_));
 sky130_fd_sc_hd__nand2_1 _05198_ (.A(net60),
    .B(net28),
    .Y(_02630_));
 sky130_fd_sc_hd__and3_1 _05199_ (.A(net60),
    .B(net28),
    .C(_02619_),
    .X(_02641_));
 sky130_fd_sc_hd__xnor2_1 _05200_ (.A(_02619_),
    .B(_02630_),
    .Y(_02652_));
 sky130_fd_sc_hd__xor2_1 _05201_ (.A(_02388_),
    .B(_02652_),
    .X(_02663_));
 sky130_fd_sc_hd__nand2_1 _05202_ (.A(net61),
    .B(net27),
    .Y(_02674_));
 sky130_fd_sc_hd__and3_1 _05203_ (.A(net61),
    .B(net27),
    .C(_02663_),
    .X(_02685_));
 sky130_fd_sc_hd__xnor2_1 _05204_ (.A(_02663_),
    .B(_02674_),
    .Y(_02696_));
 sky130_fd_sc_hd__xor2_1 _05205_ (.A(_02377_),
    .B(_02696_),
    .X(_02707_));
 sky130_fd_sc_hd__nand2_1 _05206_ (.A(net26),
    .B(net62),
    .Y(_02718_));
 sky130_fd_sc_hd__and3_1 _05207_ (.A(net26),
    .B(net62),
    .C(_02707_),
    .X(_02729_));
 sky130_fd_sc_hd__xnor2_1 _05208_ (.A(_02707_),
    .B(_02718_),
    .Y(_02740_));
 sky130_fd_sc_hd__xor2_1 _05209_ (.A(_02366_),
    .B(_02740_),
    .X(_02751_));
 sky130_fd_sc_hd__nand2_1 _05210_ (.A(net23),
    .B(net63),
    .Y(_02762_));
 sky130_fd_sc_hd__and3_1 _05211_ (.A(net23),
    .B(net63),
    .C(_02751_),
    .X(_02773_));
 sky130_fd_sc_hd__xnor2_1 _05212_ (.A(_02751_),
    .B(_02762_),
    .Y(_02784_));
 sky130_fd_sc_hd__xor2_1 _05213_ (.A(_02355_),
    .B(_02784_),
    .X(_02795_));
 sky130_fd_sc_hd__nand2_1 _05214_ (.A(net64),
    .B(net12),
    .Y(_02806_));
 sky130_fd_sc_hd__and3_1 _05215_ (.A(net64),
    .B(net12),
    .C(_02795_),
    .X(_02817_));
 sky130_fd_sc_hd__xnor2_1 _05216_ (.A(_02795_),
    .B(_02806_),
    .Y(_02828_));
 sky130_fd_sc_hd__xor2_1 _05217_ (.A(_02344_),
    .B(_02828_),
    .X(_02839_));
 sky130_fd_sc_hd__and3_1 _05218_ (.A(net34),
    .B(net1),
    .C(_02839_),
    .X(_02850_));
 sky130_fd_sc_hd__a21o_1 _05219_ (.A1(_02344_),
    .A2(_02828_),
    .B1(_02817_),
    .X(_02861_));
 sky130_fd_sc_hd__a21o_1 _05220_ (.A1(_02355_),
    .A2(_02784_),
    .B1(_02773_),
    .X(_02872_));
 sky130_fd_sc_hd__a21o_1 _05221_ (.A1(_02366_),
    .A2(_02740_),
    .B1(_02729_),
    .X(_02883_));
 sky130_fd_sc_hd__a21o_1 _05222_ (.A1(_02377_),
    .A2(_02696_),
    .B1(_02685_),
    .X(_02894_));
 sky130_fd_sc_hd__a21o_1 _05223_ (.A1(_02388_),
    .A2(_02652_),
    .B1(_02641_),
    .X(_02905_));
 sky130_fd_sc_hd__a21o_1 _05224_ (.A1(_02399_),
    .A2(_02608_),
    .B1(_02597_),
    .X(_02916_));
 sky130_fd_sc_hd__a21o_1 _05225_ (.A1(_02410_),
    .A2(_02564_),
    .B1(_02553_),
    .X(_02927_));
 sky130_fd_sc_hd__a21o_1 _05226_ (.A1(_02421_),
    .A2(_02509_),
    .B1(_02498_),
    .X(_02938_));
 sky130_fd_sc_hd__a22o_1 _05227_ (.A1(net33),
    .A2(net3),
    .B1(net2),
    .B2(net44),
    .X(_02949_));
 sky130_fd_sc_hd__and3_1 _05228_ (.A(net44),
    .B(net3),
    .C(net2),
    .X(_02960_));
 sky130_fd_sc_hd__a21bo_1 _05229_ (.A1(net33),
    .A2(_02960_),
    .B1_N(_02949_),
    .X(_02971_));
 sky130_fd_sc_hd__a21o_1 _05230_ (.A1(_02443_),
    .A2(_02465_),
    .B1(_02432_),
    .X(_02982_));
 sky130_fd_sc_hd__xnor2_1 _05231_ (.A(_02971_),
    .B(_02982_),
    .Y(_02993_));
 sky130_fd_sc_hd__nand2_1 _05232_ (.A(net55),
    .B(net32),
    .Y(_03004_));
 sky130_fd_sc_hd__and3_1 _05233_ (.A(net55),
    .B(net32),
    .C(_02993_),
    .X(_03015_));
 sky130_fd_sc_hd__nand2b_1 _05234_ (.A_N(_02993_),
    .B(_03004_),
    .Y(_03026_));
 sky130_fd_sc_hd__xor2_1 _05235_ (.A(_02993_),
    .B(_03004_),
    .X(_03037_));
 sky130_fd_sc_hd__xnor2_1 _05236_ (.A(_02938_),
    .B(_03037_),
    .Y(_03048_));
 sky130_fd_sc_hd__nand2_1 _05237_ (.A(net58),
    .B(net31),
    .Y(_03059_));
 sky130_fd_sc_hd__and3_1 _05238_ (.A(net58),
    .B(net31),
    .C(_03048_),
    .X(_03070_));
 sky130_fd_sc_hd__xnor2_1 _05239_ (.A(_03048_),
    .B(_03059_),
    .Y(_03081_));
 sky130_fd_sc_hd__xor2_1 _05240_ (.A(_02927_),
    .B(_03081_),
    .X(_03092_));
 sky130_fd_sc_hd__nand2_1 _05241_ (.A(net59),
    .B(net30),
    .Y(_03103_));
 sky130_fd_sc_hd__and3_1 _05242_ (.A(net59),
    .B(net30),
    .C(_03092_),
    .X(_03114_));
 sky130_fd_sc_hd__xnor2_1 _05243_ (.A(_03092_),
    .B(_03103_),
    .Y(_03125_));
 sky130_fd_sc_hd__xor2_1 _05244_ (.A(_02916_),
    .B(_03125_),
    .X(_03136_));
 sky130_fd_sc_hd__nand2_1 _05245_ (.A(net60),
    .B(net29),
    .Y(_03147_));
 sky130_fd_sc_hd__and3_1 _05246_ (.A(net60),
    .B(net29),
    .C(_03136_),
    .X(_03158_));
 sky130_fd_sc_hd__xnor2_1 _05247_ (.A(_03136_),
    .B(_03147_),
    .Y(_03169_));
 sky130_fd_sc_hd__xor2_1 _05248_ (.A(_02905_),
    .B(_03169_),
    .X(_03180_));
 sky130_fd_sc_hd__nand2_1 _05249_ (.A(net61),
    .B(net28),
    .Y(_03191_));
 sky130_fd_sc_hd__and3_1 _05250_ (.A(net61),
    .B(net28),
    .C(_03180_),
    .X(_03202_));
 sky130_fd_sc_hd__xnor2_1 _05251_ (.A(_03180_),
    .B(_03191_),
    .Y(_03213_));
 sky130_fd_sc_hd__xor2_1 _05252_ (.A(_02894_),
    .B(_03213_),
    .X(_03224_));
 sky130_fd_sc_hd__nand2_1 _05253_ (.A(net62),
    .B(net27),
    .Y(_03235_));
 sky130_fd_sc_hd__and3_1 _05254_ (.A(net62),
    .B(net27),
    .C(_03224_),
    .X(_03246_));
 sky130_fd_sc_hd__xnor2_1 _05255_ (.A(_03224_),
    .B(_03235_),
    .Y(_03257_));
 sky130_fd_sc_hd__xor2_1 _05256_ (.A(_02883_),
    .B(_03257_),
    .X(_03268_));
 sky130_fd_sc_hd__nand2_1 _05257_ (.A(net26),
    .B(net63),
    .Y(_03279_));
 sky130_fd_sc_hd__and3_1 _05258_ (.A(net26),
    .B(net63),
    .C(_03268_),
    .X(_03290_));
 sky130_fd_sc_hd__xnor2_1 _05259_ (.A(_03268_),
    .B(_03279_),
    .Y(_03301_));
 sky130_fd_sc_hd__xor2_1 _05260_ (.A(_02872_),
    .B(_03301_),
    .X(_03312_));
 sky130_fd_sc_hd__nand2_1 _05261_ (.A(net64),
    .B(net23),
    .Y(_03323_));
 sky130_fd_sc_hd__and3_1 _05262_ (.A(net64),
    .B(net23),
    .C(_03312_),
    .X(_03334_));
 sky130_fd_sc_hd__xnor2_1 _05263_ (.A(_03312_),
    .B(_03323_),
    .Y(_03345_));
 sky130_fd_sc_hd__xor2_1 _05264_ (.A(_02861_),
    .B(_03345_),
    .X(_03356_));
 sky130_fd_sc_hd__nand2_1 _05265_ (.A(net34),
    .B(net12),
    .Y(_03367_));
 sky130_fd_sc_hd__and3_1 _05266_ (.A(net34),
    .B(net12),
    .C(_03356_),
    .X(_03378_));
 sky130_fd_sc_hd__xnor2_1 _05267_ (.A(_03356_),
    .B(_03367_),
    .Y(_03389_));
 sky130_fd_sc_hd__xor2_1 _05268_ (.A(_02850_),
    .B(_03389_),
    .X(_03400_));
 sky130_fd_sc_hd__and3_1 _05269_ (.A(net35),
    .B(net1),
    .C(_03400_),
    .X(_03411_));
 sky130_fd_sc_hd__a21o_1 _05270_ (.A1(_02850_),
    .A2(_03389_),
    .B1(_03378_),
    .X(_03422_));
 sky130_fd_sc_hd__a21o_1 _05271_ (.A1(_02861_),
    .A2(_03345_),
    .B1(_03334_),
    .X(_03433_));
 sky130_fd_sc_hd__a21o_1 _05272_ (.A1(_02872_),
    .A2(_03301_),
    .B1(_03290_),
    .X(_03444_));
 sky130_fd_sc_hd__nand2_1 _05273_ (.A(net63),
    .B(net27),
    .Y(_03455_));
 sky130_fd_sc_hd__a21o_1 _05274_ (.A1(_02883_),
    .A2(_03257_),
    .B1(_03246_),
    .X(_03466_));
 sky130_fd_sc_hd__nand2_1 _05275_ (.A(net62),
    .B(net28),
    .Y(_03477_));
 sky130_fd_sc_hd__a21o_1 _05276_ (.A1(_02894_),
    .A2(_03213_),
    .B1(_03202_),
    .X(_03488_));
 sky130_fd_sc_hd__nand2_1 _05277_ (.A(net61),
    .B(net29),
    .Y(_03499_));
 sky130_fd_sc_hd__a21o_1 _05278_ (.A1(_02905_),
    .A2(_03169_),
    .B1(_03158_),
    .X(_03510_));
 sky130_fd_sc_hd__nand2_1 _05279_ (.A(net60),
    .B(net30),
    .Y(_03521_));
 sky130_fd_sc_hd__a21o_1 _05280_ (.A1(_02916_),
    .A2(_03125_),
    .B1(_03114_),
    .X(_03532_));
 sky130_fd_sc_hd__nand2_1 _05281_ (.A(net59),
    .B(net31),
    .Y(_03543_));
 sky130_fd_sc_hd__a21o_1 _05282_ (.A1(_02927_),
    .A2(_03081_),
    .B1(_03070_),
    .X(_03554_));
 sky130_fd_sc_hd__nand2_1 _05283_ (.A(net58),
    .B(net32),
    .Y(_03565_));
 sky130_fd_sc_hd__a21o_1 _05284_ (.A1(_02938_),
    .A2(_03026_),
    .B1(_03015_),
    .X(_03576_));
 sky130_fd_sc_hd__nand2_1 _05285_ (.A(net55),
    .B(net2),
    .Y(_03587_));
 sky130_fd_sc_hd__a22o_1 _05286_ (.A1(net33),
    .A2(net4),
    .B1(net3),
    .B2(net44),
    .X(_03598_));
 sky130_fd_sc_hd__and3_1 _05287_ (.A(net44),
    .B(net4),
    .C(net3),
    .X(_03609_));
 sky130_fd_sc_hd__a21bo_1 _05288_ (.A1(net33),
    .A2(_03609_),
    .B1_N(_03598_),
    .X(_03620_));
 sky130_fd_sc_hd__a22o_1 _05289_ (.A1(net33),
    .A2(_02960_),
    .B1(_02982_),
    .B2(_02949_),
    .X(_03631_));
 sky130_fd_sc_hd__xnor2_1 _05290_ (.A(_03620_),
    .B(_03631_),
    .Y(_03642_));
 sky130_fd_sc_hd__and3_1 _05291_ (.A(net55),
    .B(net2),
    .C(_03642_),
    .X(_03653_));
 sky130_fd_sc_hd__xnor2_1 _05292_ (.A(_03587_),
    .B(_03642_),
    .Y(_03664_));
 sky130_fd_sc_hd__xor2_1 _05293_ (.A(_03576_),
    .B(_03664_),
    .X(_03675_));
 sky130_fd_sc_hd__and3_1 _05294_ (.A(net58),
    .B(net32),
    .C(_03675_),
    .X(_03686_));
 sky130_fd_sc_hd__xnor2_1 _05295_ (.A(_03565_),
    .B(_03675_),
    .Y(_03697_));
 sky130_fd_sc_hd__xor2_1 _05296_ (.A(_03554_),
    .B(_03697_),
    .X(_03708_));
 sky130_fd_sc_hd__and3_1 _05297_ (.A(net59),
    .B(net31),
    .C(_03708_),
    .X(_03719_));
 sky130_fd_sc_hd__xnor2_1 _05298_ (.A(_03543_),
    .B(_03708_),
    .Y(_03730_));
 sky130_fd_sc_hd__xor2_1 _05299_ (.A(_03532_),
    .B(_03730_),
    .X(_03741_));
 sky130_fd_sc_hd__and3_1 _05300_ (.A(net60),
    .B(net30),
    .C(_03741_),
    .X(_03752_));
 sky130_fd_sc_hd__xnor2_1 _05301_ (.A(_03521_),
    .B(_03741_),
    .Y(_03763_));
 sky130_fd_sc_hd__xor2_1 _05302_ (.A(_03510_),
    .B(_03763_),
    .X(_03774_));
 sky130_fd_sc_hd__and3_1 _05303_ (.A(net61),
    .B(net29),
    .C(_03774_),
    .X(_03785_));
 sky130_fd_sc_hd__xnor2_1 _05304_ (.A(_03499_),
    .B(_03774_),
    .Y(_03796_));
 sky130_fd_sc_hd__xor2_1 _05305_ (.A(_03488_),
    .B(_03796_),
    .X(_03807_));
 sky130_fd_sc_hd__and3_1 _05306_ (.A(net62),
    .B(net28),
    .C(_03807_),
    .X(_03818_));
 sky130_fd_sc_hd__xnor2_1 _05307_ (.A(_03477_),
    .B(_03807_),
    .Y(_03829_));
 sky130_fd_sc_hd__xor2_1 _05308_ (.A(_03466_),
    .B(_03829_),
    .X(_03840_));
 sky130_fd_sc_hd__and3_1 _05309_ (.A(net63),
    .B(net27),
    .C(_03840_),
    .X(_03851_));
 sky130_fd_sc_hd__xnor2_1 _05310_ (.A(_03455_),
    .B(_03840_),
    .Y(_03862_));
 sky130_fd_sc_hd__xor2_1 _05311_ (.A(_03444_),
    .B(_03862_),
    .X(_03873_));
 sky130_fd_sc_hd__nand2_1 _05312_ (.A(net26),
    .B(net64),
    .Y(_03884_));
 sky130_fd_sc_hd__and3_1 _05313_ (.A(net26),
    .B(net64),
    .C(_03873_),
    .X(_03895_));
 sky130_fd_sc_hd__xnor2_1 _05314_ (.A(_03873_),
    .B(_03884_),
    .Y(_03906_));
 sky130_fd_sc_hd__xor2_1 _05315_ (.A(_03433_),
    .B(_03906_),
    .X(_03917_));
 sky130_fd_sc_hd__nand2_1 _05316_ (.A(net34),
    .B(net23),
    .Y(_03928_));
 sky130_fd_sc_hd__and3_1 _05317_ (.A(net34),
    .B(net23),
    .C(_03917_),
    .X(_03939_));
 sky130_fd_sc_hd__nand2b_1 _05318_ (.A_N(_03917_),
    .B(_03928_),
    .Y(_03950_));
 sky130_fd_sc_hd__xor2_1 _05319_ (.A(_03917_),
    .B(_03928_),
    .X(_03961_));
 sky130_fd_sc_hd__xnor2_1 _05320_ (.A(_03422_),
    .B(_03961_),
    .Y(_03972_));
 sky130_fd_sc_hd__nand2_1 _05321_ (.A(net35),
    .B(net12),
    .Y(_03983_));
 sky130_fd_sc_hd__and3_1 _05322_ (.A(net35),
    .B(net12),
    .C(_03972_),
    .X(_03994_));
 sky130_fd_sc_hd__xnor2_1 _05323_ (.A(_03972_),
    .B(_03983_),
    .Y(_04005_));
 sky130_fd_sc_hd__xor2_1 _05324_ (.A(_03411_),
    .B(_04005_),
    .X(_04016_));
 sky130_fd_sc_hd__and3_1 _05325_ (.A(net36),
    .B(net1),
    .C(_04016_),
    .X(_04027_));
 sky130_fd_sc_hd__a21oi_1 _05326_ (.A1(net36),
    .A2(net1),
    .B1(_04016_),
    .Y(_04038_));
 sky130_fd_sc_hd__nor2_1 _05327_ (.A(_04027_),
    .B(_04038_),
    .Y(\genblk2[11].rca.ripple_adders[12].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _05328_ (.A1(_03411_),
    .A2(_04005_),
    .B1(_03994_),
    .X(_04059_));
 sky130_fd_sc_hd__a21o_1 _05329_ (.A1(_03422_),
    .A2(_03950_),
    .B1(_03939_),
    .X(_04070_));
 sky130_fd_sc_hd__a21o_1 _05330_ (.A1(_03433_),
    .A2(_03906_),
    .B1(_03895_),
    .X(_04081_));
 sky130_fd_sc_hd__a21o_1 _05331_ (.A1(_03444_),
    .A2(_03862_),
    .B1(_03851_),
    .X(_04092_));
 sky130_fd_sc_hd__a21o_1 _05332_ (.A1(_03466_),
    .A2(_03829_),
    .B1(_03818_),
    .X(_04103_));
 sky130_fd_sc_hd__a21o_1 _05333_ (.A1(_03488_),
    .A2(_03796_),
    .B1(_03785_),
    .X(_04114_));
 sky130_fd_sc_hd__a21o_1 _05334_ (.A1(_03510_),
    .A2(_03763_),
    .B1(_03752_),
    .X(_04125_));
 sky130_fd_sc_hd__a21o_1 _05335_ (.A1(_03532_),
    .A2(_03730_),
    .B1(_03719_),
    .X(_04136_));
 sky130_fd_sc_hd__a21o_1 _05336_ (.A1(_03554_),
    .A2(_03697_),
    .B1(_03686_),
    .X(_04147_));
 sky130_fd_sc_hd__a21o_1 _05337_ (.A1(_03576_),
    .A2(_03664_),
    .B1(_03653_),
    .X(_04158_));
 sky130_fd_sc_hd__a22o_1 _05338_ (.A1(net33),
    .A2(net5),
    .B1(net44),
    .B2(net4),
    .X(_04169_));
 sky130_fd_sc_hd__and3_1 _05339_ (.A(net5),
    .B(net44),
    .C(net4),
    .X(_04180_));
 sky130_fd_sc_hd__a21bo_1 _05340_ (.A1(net33),
    .A2(_04180_),
    .B1_N(_04169_),
    .X(_04191_));
 sky130_fd_sc_hd__a22o_1 _05341_ (.A1(net33),
    .A2(_03609_),
    .B1(_03631_),
    .B2(_03598_),
    .X(_04202_));
 sky130_fd_sc_hd__xnor2_1 _05342_ (.A(_04191_),
    .B(_04202_),
    .Y(_04213_));
 sky130_fd_sc_hd__nand2_1 _05343_ (.A(net55),
    .B(net3),
    .Y(_04224_));
 sky130_fd_sc_hd__and3_1 _05344_ (.A(net55),
    .B(net3),
    .C(_04213_),
    .X(_04235_));
 sky130_fd_sc_hd__nand2b_1 _05345_ (.A_N(_04213_),
    .B(_04224_),
    .Y(_04246_));
 sky130_fd_sc_hd__xor2_1 _05346_ (.A(_04213_),
    .B(_04224_),
    .X(_04257_));
 sky130_fd_sc_hd__xnor2_1 _05347_ (.A(_04158_),
    .B(_04257_),
    .Y(_04268_));
 sky130_fd_sc_hd__nand2_1 _05348_ (.A(net58),
    .B(net2),
    .Y(_04279_));
 sky130_fd_sc_hd__and3_1 _05349_ (.A(net58),
    .B(net2),
    .C(_04268_),
    .X(_04290_));
 sky130_fd_sc_hd__xnor2_1 _05350_ (.A(_04268_),
    .B(_04279_),
    .Y(_04301_));
 sky130_fd_sc_hd__xor2_1 _05351_ (.A(_04147_),
    .B(_04301_),
    .X(_04312_));
 sky130_fd_sc_hd__nand2_1 _05352_ (.A(net59),
    .B(net32),
    .Y(_04323_));
 sky130_fd_sc_hd__and3_1 _05353_ (.A(net59),
    .B(net32),
    .C(_04312_),
    .X(_04334_));
 sky130_fd_sc_hd__xnor2_1 _05354_ (.A(_04312_),
    .B(_04323_),
    .Y(_04345_));
 sky130_fd_sc_hd__xor2_1 _05355_ (.A(_04136_),
    .B(_04345_),
    .X(_04356_));
 sky130_fd_sc_hd__nand2_1 _05356_ (.A(net60),
    .B(net31),
    .Y(_04367_));
 sky130_fd_sc_hd__and3_1 _05357_ (.A(net60),
    .B(net31),
    .C(_04356_),
    .X(_04378_));
 sky130_fd_sc_hd__xnor2_1 _05358_ (.A(_04356_),
    .B(_04367_),
    .Y(_04389_));
 sky130_fd_sc_hd__xor2_1 _05359_ (.A(_04125_),
    .B(_04389_),
    .X(_04400_));
 sky130_fd_sc_hd__nand2_1 _05360_ (.A(net61),
    .B(net30),
    .Y(_04411_));
 sky130_fd_sc_hd__and3_1 _05361_ (.A(net61),
    .B(net30),
    .C(_04400_),
    .X(_04422_));
 sky130_fd_sc_hd__xnor2_1 _05362_ (.A(_04400_),
    .B(_04411_),
    .Y(_04433_));
 sky130_fd_sc_hd__xor2_1 _05363_ (.A(_04114_),
    .B(_04433_),
    .X(_04444_));
 sky130_fd_sc_hd__nand2_1 _05364_ (.A(net62),
    .B(net29),
    .Y(_04455_));
 sky130_fd_sc_hd__and3_1 _05365_ (.A(net62),
    .B(net29),
    .C(_04444_),
    .X(_04466_));
 sky130_fd_sc_hd__xnor2_1 _05366_ (.A(_04444_),
    .B(_04455_),
    .Y(_04477_));
 sky130_fd_sc_hd__xor2_1 _05367_ (.A(_04103_),
    .B(_04477_),
    .X(_04488_));
 sky130_fd_sc_hd__nand2_1 _05368_ (.A(net28),
    .B(net63),
    .Y(_04492_));
 sky130_fd_sc_hd__and3_1 _05369_ (.A(net28),
    .B(net63),
    .C(_04488_),
    .X(_04493_));
 sky130_fd_sc_hd__xnor2_1 _05370_ (.A(_04488_),
    .B(_04492_),
    .Y(_04494_));
 sky130_fd_sc_hd__xor2_1 _05371_ (.A(_04092_),
    .B(_04494_),
    .X(_04498_));
 sky130_fd_sc_hd__nand2_1 _05372_ (.A(net64),
    .B(net27),
    .Y(_04504_));
 sky130_fd_sc_hd__and3_1 _05373_ (.A(net64),
    .B(net27),
    .C(_04498_),
    .X(_04508_));
 sky130_fd_sc_hd__xnor2_1 _05374_ (.A(_04498_),
    .B(_04504_),
    .Y(_04509_));
 sky130_fd_sc_hd__xor2_1 _05375_ (.A(_04081_),
    .B(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__nand2_1 _05376_ (.A(net26),
    .B(net34),
    .Y(_04511_));
 sky130_fd_sc_hd__and3_1 _05377_ (.A(net26),
    .B(net34),
    .C(_04510_),
    .X(_04512_));
 sky130_fd_sc_hd__xnor2_1 _05378_ (.A(_04510_),
    .B(_04511_),
    .Y(_04513_));
 sky130_fd_sc_hd__xor2_1 _05379_ (.A(_04070_),
    .B(_04513_),
    .X(_04514_));
 sky130_fd_sc_hd__nand2_1 _05380_ (.A(net23),
    .B(net35),
    .Y(_04515_));
 sky130_fd_sc_hd__and3_1 _05381_ (.A(net23),
    .B(net35),
    .C(_04514_),
    .X(_04516_));
 sky130_fd_sc_hd__xnor2_1 _05382_ (.A(_04514_),
    .B(_04515_),
    .Y(_04517_));
 sky130_fd_sc_hd__xor2_1 _05383_ (.A(_04059_),
    .B(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__nand2_1 _05384_ (.A(net12),
    .B(net36),
    .Y(_04519_));
 sky130_fd_sc_hd__and3_1 _05385_ (.A(net12),
    .B(net36),
    .C(_04518_),
    .X(_04520_));
 sky130_fd_sc_hd__xnor2_1 _05386_ (.A(_04518_),
    .B(_04519_),
    .Y(_04521_));
 sky130_fd_sc_hd__xor2_1 _05387_ (.A(_04027_),
    .B(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__and3_1 _05388_ (.A(net1),
    .B(net37),
    .C(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__a21oi_1 _05389_ (.A1(net1),
    .A2(net37),
    .B1(_04522_),
    .Y(_04524_));
 sky130_fd_sc_hd__nor2_1 _05390_ (.A(_04523_),
    .B(_04524_),
    .Y(\genblk2[12].rca.ripple_adders[13].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _05391_ (.A1(_04027_),
    .A2(_04521_),
    .B1(_04520_),
    .X(_04525_));
 sky130_fd_sc_hd__a21o_1 _05392_ (.A1(_04059_),
    .A2(_04517_),
    .B1(_04516_),
    .X(_04526_));
 sky130_fd_sc_hd__a21o_1 _05393_ (.A1(_04070_),
    .A2(_04513_),
    .B1(_04512_),
    .X(_04527_));
 sky130_fd_sc_hd__a21o_1 _05394_ (.A1(_04081_),
    .A2(_04509_),
    .B1(_04508_),
    .X(_04528_));
 sky130_fd_sc_hd__a21o_1 _05395_ (.A1(_04092_),
    .A2(_04494_),
    .B1(_04493_),
    .X(_04529_));
 sky130_fd_sc_hd__a21o_1 _05396_ (.A1(_04103_),
    .A2(_04477_),
    .B1(_04466_),
    .X(_04530_));
 sky130_fd_sc_hd__a21o_1 _05397_ (.A1(_04114_),
    .A2(_04433_),
    .B1(_04422_),
    .X(_04531_));
 sky130_fd_sc_hd__a21o_1 _05398_ (.A1(_04125_),
    .A2(_04389_),
    .B1(_04378_),
    .X(_04532_));
 sky130_fd_sc_hd__a21o_1 _05399_ (.A1(_04136_),
    .A2(_04345_),
    .B1(_04334_),
    .X(_04533_));
 sky130_fd_sc_hd__a21o_1 _05400_ (.A1(_04147_),
    .A2(_04301_),
    .B1(_04290_),
    .X(_04534_));
 sky130_fd_sc_hd__a21o_1 _05401_ (.A1(_04158_),
    .A2(_04246_),
    .B1(_04235_),
    .X(_04535_));
 sky130_fd_sc_hd__a22o_1 _05402_ (.A1(net5),
    .A2(net44),
    .B1(net6),
    .B2(net33),
    .X(_04536_));
 sky130_fd_sc_hd__and3_1 _05403_ (.A(net5),
    .B(net44),
    .C(net6),
    .X(_04537_));
 sky130_fd_sc_hd__a21bo_1 _05404_ (.A1(net33),
    .A2(_04537_),
    .B1_N(_04536_),
    .X(_04538_));
 sky130_fd_sc_hd__a22o_1 _05405_ (.A1(net33),
    .A2(_04180_),
    .B1(_04202_),
    .B2(_04169_),
    .X(_04539_));
 sky130_fd_sc_hd__xnor2_1 _05406_ (.A(_04538_),
    .B(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__nand2_1 _05407_ (.A(net4),
    .B(net55),
    .Y(_04541_));
 sky130_fd_sc_hd__and3_1 _05408_ (.A(net4),
    .B(net55),
    .C(_04540_),
    .X(_04542_));
 sky130_fd_sc_hd__nand2b_1 _05409_ (.A_N(_04540_),
    .B(_04541_),
    .Y(_04543_));
 sky130_fd_sc_hd__xor2_1 _05410_ (.A(_04540_),
    .B(_04541_),
    .X(_04544_));
 sky130_fd_sc_hd__xnor2_1 _05411_ (.A(_04535_),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__nand2_1 _05412_ (.A(net3),
    .B(net58),
    .Y(_04546_));
 sky130_fd_sc_hd__and3_1 _05413_ (.A(net3),
    .B(net58),
    .C(_04545_),
    .X(_04547_));
 sky130_fd_sc_hd__xnor2_1 _05414_ (.A(_04545_),
    .B(_04546_),
    .Y(_04548_));
 sky130_fd_sc_hd__xor2_1 _05415_ (.A(_04534_),
    .B(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__nand2_1 _05416_ (.A(net2),
    .B(net59),
    .Y(_04550_));
 sky130_fd_sc_hd__and3_1 _05417_ (.A(net2),
    .B(net59),
    .C(_04549_),
    .X(_04551_));
 sky130_fd_sc_hd__xnor2_1 _05418_ (.A(_04549_),
    .B(_04550_),
    .Y(_04552_));
 sky130_fd_sc_hd__xor2_1 _05419_ (.A(_04533_),
    .B(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__nand2_1 _05420_ (.A(net32),
    .B(net60),
    .Y(_04554_));
 sky130_fd_sc_hd__and3_1 _05421_ (.A(net32),
    .B(net60),
    .C(_04553_),
    .X(_04555_));
 sky130_fd_sc_hd__xnor2_1 _05422_ (.A(_04553_),
    .B(_04554_),
    .Y(_04556_));
 sky130_fd_sc_hd__xor2_1 _05423_ (.A(_04532_),
    .B(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__nand2_1 _05424_ (.A(net31),
    .B(net61),
    .Y(_04558_));
 sky130_fd_sc_hd__and3_1 _05425_ (.A(net31),
    .B(net61),
    .C(_04557_),
    .X(_04559_));
 sky130_fd_sc_hd__xnor2_1 _05426_ (.A(_04557_),
    .B(_04558_),
    .Y(_04560_));
 sky130_fd_sc_hd__xor2_1 _05427_ (.A(_04531_),
    .B(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__nand2_1 _05428_ (.A(net30),
    .B(net62),
    .Y(_04562_));
 sky130_fd_sc_hd__and3_1 _05429_ (.A(net30),
    .B(net62),
    .C(_04561_),
    .X(_04563_));
 sky130_fd_sc_hd__xnor2_1 _05430_ (.A(_04561_),
    .B(_04562_),
    .Y(_04564_));
 sky130_fd_sc_hd__xor2_1 _05431_ (.A(_04530_),
    .B(_04564_),
    .X(_04565_));
 sky130_fd_sc_hd__nand2_1 _05432_ (.A(net29),
    .B(net63),
    .Y(_04566_));
 sky130_fd_sc_hd__and3_1 _05433_ (.A(net29),
    .B(net63),
    .C(_04565_),
    .X(_04567_));
 sky130_fd_sc_hd__xnor2_1 _05434_ (.A(_04565_),
    .B(_04566_),
    .Y(_04568_));
 sky130_fd_sc_hd__xor2_1 _05435_ (.A(_04529_),
    .B(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__nand2_1 _05436_ (.A(net64),
    .B(net28),
    .Y(_04570_));
 sky130_fd_sc_hd__and3_1 _05437_ (.A(net64),
    .B(net28),
    .C(_04569_),
    .X(_04571_));
 sky130_fd_sc_hd__xnor2_1 _05438_ (.A(_04569_),
    .B(_04570_),
    .Y(_04572_));
 sky130_fd_sc_hd__xor2_1 _05439_ (.A(_04528_),
    .B(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__nand2_1 _05440_ (.A(net34),
    .B(net27),
    .Y(_04574_));
 sky130_fd_sc_hd__and3_1 _05441_ (.A(net34),
    .B(net27),
    .C(_04573_),
    .X(_04575_));
 sky130_fd_sc_hd__xnor2_1 _05442_ (.A(_04573_),
    .B(_04574_),
    .Y(_04576_));
 sky130_fd_sc_hd__xor2_1 _05443_ (.A(_04527_),
    .B(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__nand2_1 _05444_ (.A(net26),
    .B(net35),
    .Y(_04578_));
 sky130_fd_sc_hd__and3_1 _05445_ (.A(net26),
    .B(net35),
    .C(_04577_),
    .X(_04579_));
 sky130_fd_sc_hd__xnor2_1 _05446_ (.A(_04577_),
    .B(_04578_),
    .Y(_04580_));
 sky130_fd_sc_hd__xnor2_1 _05447_ (.A(_04526_),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__nand2_1 _05448_ (.A(net23),
    .B(net36),
    .Y(_04582_));
 sky130_fd_sc_hd__nor2_1 _05449_ (.A(_04581_),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__xor2_1 _05450_ (.A(_04581_),
    .B(_04582_),
    .X(_04584_));
 sky130_fd_sc_hd__xnor2_1 _05451_ (.A(_04525_),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__nand2_1 _05452_ (.A(net12),
    .B(net37),
    .Y(_04586_));
 sky130_fd_sc_hd__nor2_1 _05453_ (.A(_04585_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__xor2_1 _05454_ (.A(_04585_),
    .B(_04586_),
    .X(_04588_));
 sky130_fd_sc_hd__xor2_1 _05455_ (.A(_04523_),
    .B(_04588_),
    .X(_04589_));
 sky130_fd_sc_hd__and3_1 _05456_ (.A(net1),
    .B(net38),
    .C(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__a21oi_1 _05457_ (.A1(net1),
    .A2(net38),
    .B1(_04589_),
    .Y(_04591_));
 sky130_fd_sc_hd__nor2_1 _05458_ (.A(_04590_),
    .B(_04591_),
    .Y(\genblk2[13].rca.ripple_adders[14].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _05459_ (.A1(_04523_),
    .A2(_04588_),
    .B1(_04587_),
    .X(_04592_));
 sky130_fd_sc_hd__a21o_1 _05460_ (.A1(_04525_),
    .A2(_04584_),
    .B1(_04583_),
    .X(_04593_));
 sky130_fd_sc_hd__a21o_1 _05461_ (.A1(_04526_),
    .A2(_04580_),
    .B1(_04579_),
    .X(_04594_));
 sky130_fd_sc_hd__a21o_1 _05462_ (.A1(_04527_),
    .A2(_04576_),
    .B1(_04575_),
    .X(_04595_));
 sky130_fd_sc_hd__a21o_1 _05463_ (.A1(_04528_),
    .A2(_04572_),
    .B1(_04571_),
    .X(_04596_));
 sky130_fd_sc_hd__a21o_1 _05464_ (.A1(_04529_),
    .A2(_04568_),
    .B1(_04567_),
    .X(_04597_));
 sky130_fd_sc_hd__a21o_1 _05465_ (.A1(_04530_),
    .A2(_04564_),
    .B1(_04563_),
    .X(_04598_));
 sky130_fd_sc_hd__a21o_1 _05466_ (.A1(_04531_),
    .A2(_04560_),
    .B1(_04559_),
    .X(_04599_));
 sky130_fd_sc_hd__a21o_1 _05467_ (.A1(_04532_),
    .A2(_04556_),
    .B1(_04555_),
    .X(_04600_));
 sky130_fd_sc_hd__a21o_1 _05468_ (.A1(_04533_),
    .A2(_04552_),
    .B1(_04551_),
    .X(_04601_));
 sky130_fd_sc_hd__a21o_1 _05469_ (.A1(_04534_),
    .A2(_04548_),
    .B1(_04547_),
    .X(_04602_));
 sky130_fd_sc_hd__a21o_1 _05470_ (.A1(_04535_),
    .A2(_04543_),
    .B1(_04542_),
    .X(_04603_));
 sky130_fd_sc_hd__a22o_1 _05471_ (.A1(net44),
    .A2(net6),
    .B1(net7),
    .B2(net33),
    .X(_04604_));
 sky130_fd_sc_hd__and3_1 _05472_ (.A(net44),
    .B(net6),
    .C(net7),
    .X(_04605_));
 sky130_fd_sc_hd__a21bo_1 _05473_ (.A1(net33),
    .A2(_04605_),
    .B1_N(_04604_),
    .X(_04606_));
 sky130_fd_sc_hd__a22o_1 _05474_ (.A1(net33),
    .A2(_04537_),
    .B1(_04539_),
    .B2(_04536_),
    .X(_04607_));
 sky130_fd_sc_hd__xnor2_1 _05475_ (.A(_04606_),
    .B(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__nand2_1 _05476_ (.A(net5),
    .B(net55),
    .Y(_04609_));
 sky130_fd_sc_hd__and3_1 _05477_ (.A(net5),
    .B(net55),
    .C(_04608_),
    .X(_04610_));
 sky130_fd_sc_hd__nand2b_1 _05478_ (.A_N(_04608_),
    .B(_04609_),
    .Y(_04611_));
 sky130_fd_sc_hd__xor2_1 _05479_ (.A(_04608_),
    .B(_04609_),
    .X(_04612_));
 sky130_fd_sc_hd__xnor2_1 _05480_ (.A(_04603_),
    .B(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__nand2_1 _05481_ (.A(net4),
    .B(net58),
    .Y(_04614_));
 sky130_fd_sc_hd__and3_1 _05482_ (.A(net4),
    .B(net58),
    .C(_04613_),
    .X(_04615_));
 sky130_fd_sc_hd__xnor2_1 _05483_ (.A(_04613_),
    .B(_04614_),
    .Y(_04616_));
 sky130_fd_sc_hd__xor2_1 _05484_ (.A(_04602_),
    .B(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__nand2_1 _05485_ (.A(net3),
    .B(net59),
    .Y(_04618_));
 sky130_fd_sc_hd__and3_1 _05486_ (.A(net3),
    .B(net59),
    .C(_04617_),
    .X(_04619_));
 sky130_fd_sc_hd__xnor2_1 _05487_ (.A(_04617_),
    .B(_04618_),
    .Y(_04620_));
 sky130_fd_sc_hd__xor2_1 _05488_ (.A(_04601_),
    .B(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__nand2_1 _05489_ (.A(net2),
    .B(net60),
    .Y(_04622_));
 sky130_fd_sc_hd__and3_1 _05490_ (.A(net2),
    .B(net60),
    .C(_04621_),
    .X(_04623_));
 sky130_fd_sc_hd__xnor2_1 _05491_ (.A(_04621_),
    .B(_04622_),
    .Y(_04624_));
 sky130_fd_sc_hd__xor2_1 _05492_ (.A(_04600_),
    .B(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__nand2_1 _05493_ (.A(net32),
    .B(net61),
    .Y(_04626_));
 sky130_fd_sc_hd__and3_1 _05494_ (.A(net32),
    .B(net61),
    .C(_04625_),
    .X(_04627_));
 sky130_fd_sc_hd__xnor2_1 _05495_ (.A(_04625_),
    .B(_04626_),
    .Y(_04628_));
 sky130_fd_sc_hd__xor2_1 _05496_ (.A(_04599_),
    .B(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__nand2_1 _05497_ (.A(net31),
    .B(net62),
    .Y(_04630_));
 sky130_fd_sc_hd__and3_1 _05498_ (.A(net31),
    .B(net62),
    .C(_04629_),
    .X(_04631_));
 sky130_fd_sc_hd__xnor2_1 _05499_ (.A(_04629_),
    .B(_04630_),
    .Y(_04632_));
 sky130_fd_sc_hd__xor2_1 _05500_ (.A(_04598_),
    .B(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__nand2_1 _05501_ (.A(net30),
    .B(net63),
    .Y(_04634_));
 sky130_fd_sc_hd__and3_1 _05502_ (.A(net30),
    .B(net63),
    .C(_04633_),
    .X(_04635_));
 sky130_fd_sc_hd__xnor2_1 _05503_ (.A(_04633_),
    .B(_04634_),
    .Y(_04636_));
 sky130_fd_sc_hd__xor2_1 _05504_ (.A(_04597_),
    .B(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__nand2_1 _05505_ (.A(net64),
    .B(net29),
    .Y(_04638_));
 sky130_fd_sc_hd__and3_1 _05506_ (.A(net64),
    .B(net29),
    .C(_04637_),
    .X(_04639_));
 sky130_fd_sc_hd__xnor2_1 _05507_ (.A(_04637_),
    .B(_04638_),
    .Y(_04640_));
 sky130_fd_sc_hd__xor2_1 _05508_ (.A(_04596_),
    .B(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__nand2_1 _05509_ (.A(net34),
    .B(net28),
    .Y(_04642_));
 sky130_fd_sc_hd__and3_1 _05510_ (.A(net34),
    .B(net28),
    .C(_04641_),
    .X(_04643_));
 sky130_fd_sc_hd__xnor2_1 _05511_ (.A(_04641_),
    .B(_04642_),
    .Y(_04644_));
 sky130_fd_sc_hd__xnor2_1 _05512_ (.A(_04595_),
    .B(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__nand2_1 _05513_ (.A(net35),
    .B(net27),
    .Y(_04646_));
 sky130_fd_sc_hd__nor2_1 _05514_ (.A(_04645_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__xor2_1 _05515_ (.A(_04645_),
    .B(_04646_),
    .X(_04648_));
 sky130_fd_sc_hd__xnor2_1 _05516_ (.A(_04594_),
    .B(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_1 _05517_ (.A(net26),
    .B(net36),
    .Y(_04650_));
 sky130_fd_sc_hd__nor2_1 _05518_ (.A(_04649_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__xor2_1 _05519_ (.A(_04649_),
    .B(_04650_),
    .X(_04652_));
 sky130_fd_sc_hd__xnor2_1 _05520_ (.A(_04593_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__nand2_1 _05521_ (.A(net23),
    .B(net37),
    .Y(_04654_));
 sky130_fd_sc_hd__nor2_1 _05522_ (.A(_04653_),
    .B(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__xor2_1 _05523_ (.A(_04653_),
    .B(_04654_),
    .X(_04656_));
 sky130_fd_sc_hd__xnor2_1 _05524_ (.A(_04592_),
    .B(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__nand2_1 _05525_ (.A(net12),
    .B(net38),
    .Y(_04658_));
 sky130_fd_sc_hd__nor2_1 _05526_ (.A(_04657_),
    .B(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__xor2_1 _05527_ (.A(_04657_),
    .B(_04658_),
    .X(_04660_));
 sky130_fd_sc_hd__xor2_1 _05528_ (.A(_04590_),
    .B(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__and3_1 _05529_ (.A(net1),
    .B(net39),
    .C(_04661_),
    .X(_04662_));
 sky130_fd_sc_hd__a21oi_1 _05530_ (.A1(net1),
    .A2(net39),
    .B1(_04661_),
    .Y(_04663_));
 sky130_fd_sc_hd__nor2_1 _05531_ (.A(_04662_),
    .B(_04663_),
    .Y(\genblk2[14].rca.ripple_adders[15].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _05532_ (.A1(_04590_),
    .A2(_04660_),
    .B1(_04659_),
    .X(_04664_));
 sky130_fd_sc_hd__a21o_1 _05533_ (.A1(_04592_),
    .A2(_04656_),
    .B1(_04655_),
    .X(_04665_));
 sky130_fd_sc_hd__a21o_1 _05534_ (.A1(_04593_),
    .A2(_04652_),
    .B1(_04651_),
    .X(_04666_));
 sky130_fd_sc_hd__a21o_1 _05535_ (.A1(_04594_),
    .A2(_04648_),
    .B1(_04647_),
    .X(_04667_));
 sky130_fd_sc_hd__a21o_1 _05536_ (.A1(_04595_),
    .A2(_04644_),
    .B1(_04643_),
    .X(_04668_));
 sky130_fd_sc_hd__a21o_1 _05537_ (.A1(_04596_),
    .A2(_04640_),
    .B1(_04639_),
    .X(_04669_));
 sky130_fd_sc_hd__a21o_1 _05538_ (.A1(_04597_),
    .A2(_04636_),
    .B1(_04635_),
    .X(_04670_));
 sky130_fd_sc_hd__a21o_1 _05539_ (.A1(_04598_),
    .A2(_04632_),
    .B1(_04631_),
    .X(_04671_));
 sky130_fd_sc_hd__a21o_1 _05540_ (.A1(_04599_),
    .A2(_04628_),
    .B1(_04627_),
    .X(_04672_));
 sky130_fd_sc_hd__a21o_1 _05541_ (.A1(_04600_),
    .A2(_04624_),
    .B1(_04623_),
    .X(_04673_));
 sky130_fd_sc_hd__a21o_1 _05542_ (.A1(_04601_),
    .A2(_04620_),
    .B1(_04619_),
    .X(_04674_));
 sky130_fd_sc_hd__a21o_1 _05543_ (.A1(_04602_),
    .A2(_04616_),
    .B1(_04615_),
    .X(_04675_));
 sky130_fd_sc_hd__a21o_1 _05544_ (.A1(_04603_),
    .A2(_04611_),
    .B1(_04610_),
    .X(_04676_));
 sky130_fd_sc_hd__a22o_1 _05545_ (.A1(net44),
    .A2(net7),
    .B1(net8),
    .B2(net33),
    .X(_04677_));
 sky130_fd_sc_hd__and3_1 _05546_ (.A(net44),
    .B(net7),
    .C(net8),
    .X(_04678_));
 sky130_fd_sc_hd__a21bo_1 _05547_ (.A1(net33),
    .A2(_04678_),
    .B1_N(_04677_),
    .X(_04679_));
 sky130_fd_sc_hd__a22o_1 _05548_ (.A1(net33),
    .A2(_04605_),
    .B1(_04607_),
    .B2(_04604_),
    .X(_04680_));
 sky130_fd_sc_hd__xnor2_1 _05549_ (.A(_04679_),
    .B(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__nand2_1 _05550_ (.A(net55),
    .B(net6),
    .Y(_04682_));
 sky130_fd_sc_hd__and3_1 _05551_ (.A(net55),
    .B(net6),
    .C(_04681_),
    .X(_04683_));
 sky130_fd_sc_hd__nand2b_1 _05552_ (.A_N(_04681_),
    .B(_04682_),
    .Y(_04684_));
 sky130_fd_sc_hd__xor2_1 _05553_ (.A(_04681_),
    .B(_04682_),
    .X(_04685_));
 sky130_fd_sc_hd__xnor2_1 _05554_ (.A(_04676_),
    .B(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__nand2_1 _05555_ (.A(net5),
    .B(net58),
    .Y(_04687_));
 sky130_fd_sc_hd__and3_1 _05556_ (.A(net5),
    .B(net58),
    .C(_04686_),
    .X(_04688_));
 sky130_fd_sc_hd__xnor2_1 _05557_ (.A(_04686_),
    .B(_04687_),
    .Y(_04689_));
 sky130_fd_sc_hd__xor2_1 _05558_ (.A(_04675_),
    .B(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__nand2_1 _05559_ (.A(net4),
    .B(net59),
    .Y(_04691_));
 sky130_fd_sc_hd__and3_1 _05560_ (.A(net4),
    .B(net59),
    .C(_04690_),
    .X(_04692_));
 sky130_fd_sc_hd__xnor2_1 _05561_ (.A(_04690_),
    .B(_04691_),
    .Y(_04693_));
 sky130_fd_sc_hd__xor2_1 _05562_ (.A(_04674_),
    .B(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__nand2_1 _05563_ (.A(net3),
    .B(net60),
    .Y(_04695_));
 sky130_fd_sc_hd__and3_1 _05564_ (.A(net3),
    .B(net60),
    .C(_04694_),
    .X(_04696_));
 sky130_fd_sc_hd__xnor2_1 _05565_ (.A(_04694_),
    .B(_04695_),
    .Y(_04697_));
 sky130_fd_sc_hd__xor2_1 _05566_ (.A(_04673_),
    .B(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__nand2_1 _05567_ (.A(net2),
    .B(net61),
    .Y(_04699_));
 sky130_fd_sc_hd__and3_1 _05568_ (.A(net2),
    .B(net61),
    .C(_04698_),
    .X(_04700_));
 sky130_fd_sc_hd__xnor2_1 _05569_ (.A(_04698_),
    .B(_04699_),
    .Y(_04701_));
 sky130_fd_sc_hd__xor2_1 _05570_ (.A(_04672_),
    .B(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__nand2_1 _05571_ (.A(net32),
    .B(net62),
    .Y(_04703_));
 sky130_fd_sc_hd__and3_1 _05572_ (.A(net32),
    .B(net62),
    .C(_04702_),
    .X(_04704_));
 sky130_fd_sc_hd__xnor2_1 _05573_ (.A(_04702_),
    .B(_04703_),
    .Y(_04705_));
 sky130_fd_sc_hd__xor2_1 _05574_ (.A(_04671_),
    .B(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__nand2_1 _05575_ (.A(net31),
    .B(net63),
    .Y(_04707_));
 sky130_fd_sc_hd__and3_1 _05576_ (.A(net31),
    .B(net63),
    .C(_04706_),
    .X(_04708_));
 sky130_fd_sc_hd__xnor2_1 _05577_ (.A(_04706_),
    .B(_04707_),
    .Y(_04709_));
 sky130_fd_sc_hd__xor2_1 _05578_ (.A(_04670_),
    .B(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__nand2_1 _05579_ (.A(net64),
    .B(net30),
    .Y(_04711_));
 sky130_fd_sc_hd__and3_1 _05580_ (.A(net64),
    .B(net30),
    .C(_04710_),
    .X(_04712_));
 sky130_fd_sc_hd__xnor2_1 _05581_ (.A(_04710_),
    .B(_04711_),
    .Y(_04713_));
 sky130_fd_sc_hd__xnor2_1 _05582_ (.A(_04669_),
    .B(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__nand2_1 _05583_ (.A(net34),
    .B(net29),
    .Y(_04715_));
 sky130_fd_sc_hd__nor2_1 _05584_ (.A(_04714_),
    .B(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__xor2_1 _05585_ (.A(_04714_),
    .B(_04715_),
    .X(_04717_));
 sky130_fd_sc_hd__xnor2_1 _05586_ (.A(_04668_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__nand2_1 _05587_ (.A(net35),
    .B(net28),
    .Y(_04719_));
 sky130_fd_sc_hd__nor2_1 _05588_ (.A(_04718_),
    .B(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__xor2_1 _05589_ (.A(_04718_),
    .B(_04719_),
    .X(_04721_));
 sky130_fd_sc_hd__xnor2_1 _05590_ (.A(_04667_),
    .B(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__nand2_1 _05591_ (.A(net36),
    .B(net27),
    .Y(_04723_));
 sky130_fd_sc_hd__nor2_1 _05592_ (.A(_04722_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__xor2_1 _05593_ (.A(_04722_),
    .B(_04723_),
    .X(_04725_));
 sky130_fd_sc_hd__xnor2_1 _05594_ (.A(_04666_),
    .B(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__nand2_1 _05595_ (.A(net26),
    .B(net37),
    .Y(_04727_));
 sky130_fd_sc_hd__nor2_1 _05596_ (.A(_04726_),
    .B(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hd__xor2_1 _05597_ (.A(_04726_),
    .B(_04727_),
    .X(_04729_));
 sky130_fd_sc_hd__xnor2_1 _05598_ (.A(_04665_),
    .B(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__nand2_1 _05599_ (.A(net23),
    .B(net38),
    .Y(_04731_));
 sky130_fd_sc_hd__nor2_1 _05600_ (.A(_04730_),
    .B(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__xor2_1 _05601_ (.A(_04730_),
    .B(_04731_),
    .X(_04733_));
 sky130_fd_sc_hd__xnor2_1 _05602_ (.A(_04664_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__nand2_1 _05603_ (.A(net12),
    .B(net39),
    .Y(_04735_));
 sky130_fd_sc_hd__nor2_1 _05604_ (.A(_04734_),
    .B(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__xor2_1 _05605_ (.A(_04734_),
    .B(_04735_),
    .X(_04737_));
 sky130_fd_sc_hd__xor2_1 _05606_ (.A(_04662_),
    .B(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__and3_1 _05607_ (.A(net1),
    .B(net40),
    .C(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__a21oi_1 _05608_ (.A1(net1),
    .A2(net40),
    .B1(_04738_),
    .Y(_04740_));
 sky130_fd_sc_hd__nor2_1 _05609_ (.A(_04739_),
    .B(_04740_),
    .Y(\genblk2[15].rca.ripple_adders[16].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _05610_ (.A1(_04662_),
    .A2(_04737_),
    .B1(_04736_),
    .X(_04741_));
 sky130_fd_sc_hd__a21o_1 _05611_ (.A1(_04664_),
    .A2(_04733_),
    .B1(_04732_),
    .X(_04742_));
 sky130_fd_sc_hd__a21o_1 _05612_ (.A1(_04665_),
    .A2(_04729_),
    .B1(_04728_),
    .X(_04743_));
 sky130_fd_sc_hd__a21o_1 _05613_ (.A1(_04666_),
    .A2(_04725_),
    .B1(_04724_),
    .X(_04744_));
 sky130_fd_sc_hd__a21o_1 _05614_ (.A1(_04667_),
    .A2(_04721_),
    .B1(_04720_),
    .X(_04745_));
 sky130_fd_sc_hd__a21o_1 _05615_ (.A1(_04668_),
    .A2(_04717_),
    .B1(_04716_),
    .X(_04746_));
 sky130_fd_sc_hd__a21o_1 _05616_ (.A1(_04669_),
    .A2(_04713_),
    .B1(_04712_),
    .X(_04747_));
 sky130_fd_sc_hd__a21o_1 _05617_ (.A1(_04670_),
    .A2(_04709_),
    .B1(_04708_),
    .X(_04748_));
 sky130_fd_sc_hd__a21o_1 _05618_ (.A1(_04671_),
    .A2(_04705_),
    .B1(_04704_),
    .X(_04749_));
 sky130_fd_sc_hd__a21o_1 _05619_ (.A1(_04672_),
    .A2(_04701_),
    .B1(_04700_),
    .X(_04750_));
 sky130_fd_sc_hd__a21o_1 _05620_ (.A1(_04673_),
    .A2(_04697_),
    .B1(_04696_),
    .X(_04751_));
 sky130_fd_sc_hd__a21o_1 _05621_ (.A1(_04674_),
    .A2(_04693_),
    .B1(_04692_),
    .X(_04752_));
 sky130_fd_sc_hd__a21o_1 _05622_ (.A1(_04675_),
    .A2(_04689_),
    .B1(_04688_),
    .X(_04753_));
 sky130_fd_sc_hd__a21o_1 _05623_ (.A1(_04676_),
    .A2(_04684_),
    .B1(_04683_),
    .X(_04754_));
 sky130_fd_sc_hd__a22o_1 _05624_ (.A1(net44),
    .A2(net8),
    .B1(net9),
    .B2(net33),
    .X(_04755_));
 sky130_fd_sc_hd__and3_1 _05625_ (.A(net44),
    .B(net8),
    .C(net9),
    .X(_04756_));
 sky130_fd_sc_hd__a21bo_1 _05626_ (.A1(net33),
    .A2(_04756_),
    .B1_N(_04755_),
    .X(_04757_));
 sky130_fd_sc_hd__a22o_1 _05627_ (.A1(net33),
    .A2(_04678_),
    .B1(_04680_),
    .B2(_04677_),
    .X(_04758_));
 sky130_fd_sc_hd__xnor2_1 _05628_ (.A(_04757_),
    .B(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__nand2_1 _05629_ (.A(net55),
    .B(net7),
    .Y(_04760_));
 sky130_fd_sc_hd__and3_1 _05630_ (.A(net55),
    .B(net7),
    .C(_04759_),
    .X(_04761_));
 sky130_fd_sc_hd__nand2b_1 _05631_ (.A_N(_04759_),
    .B(_04760_),
    .Y(_04762_));
 sky130_fd_sc_hd__xor2_1 _05632_ (.A(_04759_),
    .B(_04760_),
    .X(_04763_));
 sky130_fd_sc_hd__xnor2_1 _05633_ (.A(_04754_),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__nand2_1 _05634_ (.A(net58),
    .B(net6),
    .Y(_04765_));
 sky130_fd_sc_hd__and3_1 _05635_ (.A(net58),
    .B(net6),
    .C(_04764_),
    .X(_04766_));
 sky130_fd_sc_hd__xnor2_1 _05636_ (.A(_04764_),
    .B(_04765_),
    .Y(_04767_));
 sky130_fd_sc_hd__xor2_1 _05637_ (.A(_04753_),
    .B(_04767_),
    .X(_04768_));
 sky130_fd_sc_hd__nand2_1 _05638_ (.A(net5),
    .B(net59),
    .Y(_04769_));
 sky130_fd_sc_hd__and3_1 _05639_ (.A(net5),
    .B(net59),
    .C(_04768_),
    .X(_04770_));
 sky130_fd_sc_hd__xnor2_1 _05640_ (.A(_04768_),
    .B(_04769_),
    .Y(_04771_));
 sky130_fd_sc_hd__xor2_1 _05641_ (.A(_04752_),
    .B(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__nand2_1 _05642_ (.A(net4),
    .B(net60),
    .Y(_04773_));
 sky130_fd_sc_hd__and3_1 _05643_ (.A(net4),
    .B(net60),
    .C(_04772_),
    .X(_04774_));
 sky130_fd_sc_hd__xnor2_1 _05644_ (.A(_04772_),
    .B(_04773_),
    .Y(_04775_));
 sky130_fd_sc_hd__xor2_1 _05645_ (.A(_04751_),
    .B(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__nand2_1 _05646_ (.A(net3),
    .B(net61),
    .Y(_04777_));
 sky130_fd_sc_hd__and3_1 _05647_ (.A(net3),
    .B(net61),
    .C(_04776_),
    .X(_04778_));
 sky130_fd_sc_hd__xnor2_1 _05648_ (.A(_04776_),
    .B(_04777_),
    .Y(_04779_));
 sky130_fd_sc_hd__xor2_1 _05649_ (.A(_04750_),
    .B(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__nand2_1 _05650_ (.A(net2),
    .B(net62),
    .Y(_04781_));
 sky130_fd_sc_hd__and3_1 _05651_ (.A(net2),
    .B(net62),
    .C(_04780_),
    .X(_04782_));
 sky130_fd_sc_hd__xnor2_1 _05652_ (.A(_04780_),
    .B(_04781_),
    .Y(_04783_));
 sky130_fd_sc_hd__xor2_1 _05653_ (.A(_04749_),
    .B(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__nand2_1 _05654_ (.A(net32),
    .B(net63),
    .Y(_04785_));
 sky130_fd_sc_hd__and3_1 _05655_ (.A(net32),
    .B(net63),
    .C(_04784_),
    .X(_04786_));
 sky130_fd_sc_hd__xnor2_1 _05656_ (.A(_04784_),
    .B(_04785_),
    .Y(_04787_));
 sky130_fd_sc_hd__xor2_1 _05657_ (.A(_04748_),
    .B(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__nand2_1 _05658_ (.A(net64),
    .B(net31),
    .Y(_04789_));
 sky130_fd_sc_hd__and3_1 _05659_ (.A(net64),
    .B(net31),
    .C(_04788_),
    .X(_04790_));
 sky130_fd_sc_hd__xnor2_1 _05660_ (.A(_04788_),
    .B(_04789_),
    .Y(_04791_));
 sky130_fd_sc_hd__xnor2_1 _05661_ (.A(_04747_),
    .B(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__nand2_1 _05662_ (.A(net34),
    .B(net30),
    .Y(_04793_));
 sky130_fd_sc_hd__nor2_1 _05663_ (.A(_04792_),
    .B(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__xor2_1 _05664_ (.A(_04792_),
    .B(_04793_),
    .X(_04795_));
 sky130_fd_sc_hd__xnor2_1 _05665_ (.A(_04746_),
    .B(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__nand2_1 _05666_ (.A(net35),
    .B(net29),
    .Y(_04797_));
 sky130_fd_sc_hd__nor2_1 _05667_ (.A(_04796_),
    .B(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__xor2_1 _05668_ (.A(_04796_),
    .B(_04797_),
    .X(_04799_));
 sky130_fd_sc_hd__xnor2_1 _05669_ (.A(_04745_),
    .B(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__nand2_1 _05670_ (.A(net36),
    .B(net28),
    .Y(_04801_));
 sky130_fd_sc_hd__nor2_1 _05671_ (.A(_04800_),
    .B(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__xor2_1 _05672_ (.A(_04800_),
    .B(_04801_),
    .X(_04803_));
 sky130_fd_sc_hd__xnor2_1 _05673_ (.A(_04744_),
    .B(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__nand2_1 _05674_ (.A(net27),
    .B(net37),
    .Y(_04805_));
 sky130_fd_sc_hd__nor2_1 _05675_ (.A(_04804_),
    .B(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__xor2_1 _05676_ (.A(_04804_),
    .B(_04805_),
    .X(_04807_));
 sky130_fd_sc_hd__xnor2_1 _05677_ (.A(_04743_),
    .B(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hd__nand2_1 _05678_ (.A(net26),
    .B(net38),
    .Y(_04809_));
 sky130_fd_sc_hd__nor2_1 _05679_ (.A(_04808_),
    .B(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__xor2_1 _05680_ (.A(_04808_),
    .B(_04809_),
    .X(_04811_));
 sky130_fd_sc_hd__xnor2_1 _05681_ (.A(_04742_),
    .B(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__nand2_1 _05682_ (.A(net23),
    .B(net39),
    .Y(_04813_));
 sky130_fd_sc_hd__nor2_1 _05683_ (.A(_04812_),
    .B(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__xor2_1 _05684_ (.A(_04812_),
    .B(_04813_),
    .X(_04815_));
 sky130_fd_sc_hd__xnor2_1 _05685_ (.A(_04741_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2_1 _05686_ (.A(net12),
    .B(net40),
    .Y(_04817_));
 sky130_fd_sc_hd__nor2_1 _05687_ (.A(_04816_),
    .B(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__xor2_1 _05688_ (.A(_04816_),
    .B(_04817_),
    .X(_04819_));
 sky130_fd_sc_hd__xor2_1 _05689_ (.A(_04739_),
    .B(_04819_),
    .X(_04820_));
 sky130_fd_sc_hd__and3_1 _05690_ (.A(net1),
    .B(net41),
    .C(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__a21oi_1 _05691_ (.A1(net1),
    .A2(net41),
    .B1(_04820_),
    .Y(_04822_));
 sky130_fd_sc_hd__nor2_1 _05692_ (.A(_04821_),
    .B(_04822_),
    .Y(\genblk2[16].rca.ripple_adders[17].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _05693_ (.A1(_04739_),
    .A2(_04819_),
    .B1(_04818_),
    .X(_04823_));
 sky130_fd_sc_hd__a21o_1 _05694_ (.A1(_04741_),
    .A2(_04815_),
    .B1(_04814_),
    .X(_04824_));
 sky130_fd_sc_hd__a21o_1 _05695_ (.A1(_04742_),
    .A2(_04811_),
    .B1(_04810_),
    .X(_04825_));
 sky130_fd_sc_hd__a21o_1 _05696_ (.A1(_04743_),
    .A2(_04807_),
    .B1(_04806_),
    .X(_04826_));
 sky130_fd_sc_hd__a21o_1 _05697_ (.A1(_04744_),
    .A2(_04803_),
    .B1(_04802_),
    .X(_04827_));
 sky130_fd_sc_hd__a21o_1 _05698_ (.A1(_04745_),
    .A2(_04799_),
    .B1(_04798_),
    .X(_04828_));
 sky130_fd_sc_hd__a21o_1 _05699_ (.A1(_04746_),
    .A2(_04795_),
    .B1(_04794_),
    .X(_04829_));
 sky130_fd_sc_hd__a21o_1 _05700_ (.A1(_04747_),
    .A2(_04791_),
    .B1(_04790_),
    .X(_04830_));
 sky130_fd_sc_hd__a21o_1 _05701_ (.A1(_04748_),
    .A2(_04787_),
    .B1(_04786_),
    .X(_04831_));
 sky130_fd_sc_hd__a21o_1 _05702_ (.A1(_04749_),
    .A2(_04783_),
    .B1(_04782_),
    .X(_04832_));
 sky130_fd_sc_hd__a21o_1 _05703_ (.A1(_04750_),
    .A2(_04779_),
    .B1(_04778_),
    .X(_04833_));
 sky130_fd_sc_hd__a21o_1 _05704_ (.A1(_04751_),
    .A2(_04775_),
    .B1(_04774_),
    .X(_04834_));
 sky130_fd_sc_hd__a21o_1 _05705_ (.A1(_04752_),
    .A2(_04771_),
    .B1(_04770_),
    .X(_04835_));
 sky130_fd_sc_hd__a21o_1 _05706_ (.A1(_04753_),
    .A2(_04767_),
    .B1(_04766_),
    .X(_04836_));
 sky130_fd_sc_hd__a21o_1 _05707_ (.A1(_04754_),
    .A2(_04762_),
    .B1(_04761_),
    .X(_04837_));
 sky130_fd_sc_hd__a22o_1 _05708_ (.A1(net44),
    .A2(net9),
    .B1(net10),
    .B2(net33),
    .X(_04838_));
 sky130_fd_sc_hd__and3_1 _05709_ (.A(net44),
    .B(net9),
    .C(net10),
    .X(_04839_));
 sky130_fd_sc_hd__a21bo_1 _05710_ (.A1(net33),
    .A2(_04839_),
    .B1_N(_04838_),
    .X(_04840_));
 sky130_fd_sc_hd__a22o_1 _05711_ (.A1(net33),
    .A2(_04756_),
    .B1(_04758_),
    .B2(_04755_),
    .X(_04841_));
 sky130_fd_sc_hd__xnor2_1 _05712_ (.A(_04840_),
    .B(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__nand2_1 _05713_ (.A(net55),
    .B(net8),
    .Y(_04843_));
 sky130_fd_sc_hd__and3_1 _05714_ (.A(net55),
    .B(net8),
    .C(_04842_),
    .X(_04844_));
 sky130_fd_sc_hd__nand2b_1 _05715_ (.A_N(_04842_),
    .B(_04843_),
    .Y(_04845_));
 sky130_fd_sc_hd__xor2_1 _05716_ (.A(_04842_),
    .B(_04843_),
    .X(_04846_));
 sky130_fd_sc_hd__xnor2_1 _05717_ (.A(_04837_),
    .B(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_1 _05718_ (.A(net58),
    .B(net7),
    .Y(_04848_));
 sky130_fd_sc_hd__and3_1 _05719_ (.A(net58),
    .B(net7),
    .C(_04847_),
    .X(_04849_));
 sky130_fd_sc_hd__xnor2_1 _05720_ (.A(_04847_),
    .B(_04848_),
    .Y(_04850_));
 sky130_fd_sc_hd__xor2_1 _05721_ (.A(_04836_),
    .B(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__nand2_1 _05722_ (.A(net59),
    .B(net6),
    .Y(_04852_));
 sky130_fd_sc_hd__and3_1 _05723_ (.A(net59),
    .B(net6),
    .C(_04851_),
    .X(_04853_));
 sky130_fd_sc_hd__xnor2_1 _05724_ (.A(_04851_),
    .B(_04852_),
    .Y(_04854_));
 sky130_fd_sc_hd__xor2_1 _05725_ (.A(_04835_),
    .B(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__nand2_1 _05726_ (.A(net5),
    .B(net60),
    .Y(_04856_));
 sky130_fd_sc_hd__and3_1 _05727_ (.A(net5),
    .B(net60),
    .C(_04855_),
    .X(_04857_));
 sky130_fd_sc_hd__xnor2_1 _05728_ (.A(_04855_),
    .B(_04856_),
    .Y(_04858_));
 sky130_fd_sc_hd__xor2_1 _05729_ (.A(_04834_),
    .B(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__nand2_1 _05730_ (.A(net4),
    .B(net61),
    .Y(_04860_));
 sky130_fd_sc_hd__and3_1 _05731_ (.A(net4),
    .B(net61),
    .C(_04859_),
    .X(_04861_));
 sky130_fd_sc_hd__xnor2_1 _05732_ (.A(_04859_),
    .B(_04860_),
    .Y(_04862_));
 sky130_fd_sc_hd__xor2_1 _05733_ (.A(_04833_),
    .B(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__nand2_1 _05734_ (.A(net3),
    .B(net62),
    .Y(_04864_));
 sky130_fd_sc_hd__and3_1 _05735_ (.A(net3),
    .B(net62),
    .C(_04863_),
    .X(_04865_));
 sky130_fd_sc_hd__xnor2_1 _05736_ (.A(_04863_),
    .B(_04864_),
    .Y(_04866_));
 sky130_fd_sc_hd__xor2_1 _05737_ (.A(_04832_),
    .B(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__nand2_1 _05738_ (.A(net2),
    .B(net63),
    .Y(_04868_));
 sky130_fd_sc_hd__and3_1 _05739_ (.A(net2),
    .B(net63),
    .C(_04867_),
    .X(_04869_));
 sky130_fd_sc_hd__xnor2_1 _05740_ (.A(_04867_),
    .B(_04868_),
    .Y(_04870_));
 sky130_fd_sc_hd__xnor2_1 _05741_ (.A(_04831_),
    .B(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__nand2_1 _05742_ (.A(net64),
    .B(net32),
    .Y(_04872_));
 sky130_fd_sc_hd__nor2_1 _05743_ (.A(_04871_),
    .B(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__xor2_1 _05744_ (.A(_04871_),
    .B(_04872_),
    .X(_04874_));
 sky130_fd_sc_hd__xnor2_1 _05745_ (.A(_04830_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__nand2_1 _05746_ (.A(net34),
    .B(net31),
    .Y(_04876_));
 sky130_fd_sc_hd__nor2_1 _05747_ (.A(_04875_),
    .B(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__xor2_1 _05748_ (.A(_04875_),
    .B(_04876_),
    .X(_04878_));
 sky130_fd_sc_hd__xnor2_1 _05749_ (.A(_04829_),
    .B(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hd__nand2_1 _05750_ (.A(net35),
    .B(net30),
    .Y(_04880_));
 sky130_fd_sc_hd__nor2_1 _05751_ (.A(_04879_),
    .B(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__xor2_1 _05752_ (.A(_04879_),
    .B(_04880_),
    .X(_04882_));
 sky130_fd_sc_hd__xnor2_1 _05753_ (.A(_04828_),
    .B(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__nand2_1 _05754_ (.A(net36),
    .B(net29),
    .Y(_04884_));
 sky130_fd_sc_hd__nor2_1 _05755_ (.A(_04883_),
    .B(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__xor2_1 _05756_ (.A(_04883_),
    .B(_04884_),
    .X(_04886_));
 sky130_fd_sc_hd__xnor2_1 _05757_ (.A(_04827_),
    .B(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__nand2_1 _05758_ (.A(net28),
    .B(net37),
    .Y(_04888_));
 sky130_fd_sc_hd__nor2_1 _05759_ (.A(_04887_),
    .B(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__xor2_1 _05760_ (.A(_04887_),
    .B(_04888_),
    .X(_04890_));
 sky130_fd_sc_hd__xnor2_1 _05761_ (.A(_04826_),
    .B(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__nand2_1 _05762_ (.A(net27),
    .B(net38),
    .Y(_04892_));
 sky130_fd_sc_hd__nor2_1 _05763_ (.A(_04891_),
    .B(_04892_),
    .Y(_04893_));
 sky130_fd_sc_hd__xor2_1 _05764_ (.A(_04891_),
    .B(_04892_),
    .X(_04894_));
 sky130_fd_sc_hd__xnor2_1 _05765_ (.A(_04825_),
    .B(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__nand2_1 _05766_ (.A(net26),
    .B(net39),
    .Y(_04896_));
 sky130_fd_sc_hd__nor2_1 _05767_ (.A(_04895_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__xor2_1 _05768_ (.A(_04895_),
    .B(_04896_),
    .X(_04898_));
 sky130_fd_sc_hd__xnor2_1 _05769_ (.A(_04824_),
    .B(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__nand2_1 _05770_ (.A(net23),
    .B(net40),
    .Y(_04900_));
 sky130_fd_sc_hd__nor2_1 _05771_ (.A(_04899_),
    .B(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__xor2_1 _05772_ (.A(_04899_),
    .B(_04900_),
    .X(_04902_));
 sky130_fd_sc_hd__xnor2_1 _05773_ (.A(_04823_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__nand2_1 _05774_ (.A(net12),
    .B(net41),
    .Y(_04904_));
 sky130_fd_sc_hd__nor2_1 _05775_ (.A(_04903_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__xor2_1 _05776_ (.A(_04903_),
    .B(_04904_),
    .X(_04906_));
 sky130_fd_sc_hd__xor2_1 _05777_ (.A(_04821_),
    .B(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__and3_1 _05778_ (.A(net1),
    .B(net42),
    .C(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__a21oi_1 _05779_ (.A1(net1),
    .A2(net42),
    .B1(_04907_),
    .Y(_04909_));
 sky130_fd_sc_hd__nor2_1 _05780_ (.A(_04908_),
    .B(_04909_),
    .Y(\genblk2[17].rca.ripple_adders[18].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _05781_ (.A1(_04821_),
    .A2(_04906_),
    .B1(_04905_),
    .X(_04910_));
 sky130_fd_sc_hd__a21o_1 _05782_ (.A1(_04823_),
    .A2(_04902_),
    .B1(_04901_),
    .X(_04911_));
 sky130_fd_sc_hd__a21o_1 _05783_ (.A1(_04824_),
    .A2(_04898_),
    .B1(_04897_),
    .X(_04912_));
 sky130_fd_sc_hd__a21o_1 _05784_ (.A1(_04825_),
    .A2(_04894_),
    .B1(_04893_),
    .X(_04913_));
 sky130_fd_sc_hd__a21o_1 _05785_ (.A1(_04826_),
    .A2(_04890_),
    .B1(_04889_),
    .X(_04914_));
 sky130_fd_sc_hd__a21o_1 _05786_ (.A1(_04827_),
    .A2(_04886_),
    .B1(_04885_),
    .X(_04915_));
 sky130_fd_sc_hd__a21o_1 _05787_ (.A1(_04828_),
    .A2(_04882_),
    .B1(_04881_),
    .X(_04916_));
 sky130_fd_sc_hd__a21o_1 _05788_ (.A1(_04829_),
    .A2(_04878_),
    .B1(_04877_),
    .X(_04917_));
 sky130_fd_sc_hd__a21o_1 _05789_ (.A1(_04830_),
    .A2(_04874_),
    .B1(_04873_),
    .X(_04918_));
 sky130_fd_sc_hd__a21o_1 _05790_ (.A1(_04831_),
    .A2(_04870_),
    .B1(_04869_),
    .X(_04919_));
 sky130_fd_sc_hd__a21o_1 _05791_ (.A1(_04832_),
    .A2(_04866_),
    .B1(_04865_),
    .X(_04920_));
 sky130_fd_sc_hd__a21o_1 _05792_ (.A1(_04833_),
    .A2(_04862_),
    .B1(_04861_),
    .X(_04921_));
 sky130_fd_sc_hd__a21o_1 _05793_ (.A1(_04834_),
    .A2(_04858_),
    .B1(_04857_),
    .X(_04922_));
 sky130_fd_sc_hd__a21o_1 _05794_ (.A1(_04835_),
    .A2(_04854_),
    .B1(_04853_),
    .X(_04923_));
 sky130_fd_sc_hd__a21o_1 _05795_ (.A1(_04836_),
    .A2(_04850_),
    .B1(_04849_),
    .X(_04924_));
 sky130_fd_sc_hd__a21o_1 _05796_ (.A1(_04837_),
    .A2(_04845_),
    .B1(_04844_),
    .X(_04925_));
 sky130_fd_sc_hd__a22o_1 _05797_ (.A1(net44),
    .A2(net10),
    .B1(net11),
    .B2(net33),
    .X(_04926_));
 sky130_fd_sc_hd__and3_1 _05798_ (.A(net44),
    .B(net10),
    .C(net11),
    .X(_04927_));
 sky130_fd_sc_hd__a21bo_1 _05799_ (.A1(net33),
    .A2(_04927_),
    .B1_N(_04926_),
    .X(_04928_));
 sky130_fd_sc_hd__a22o_1 _05800_ (.A1(net33),
    .A2(_04839_),
    .B1(_04841_),
    .B2(_04838_),
    .X(_04929_));
 sky130_fd_sc_hd__xnor2_1 _05801_ (.A(_04928_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__nand2_1 _05802_ (.A(net55),
    .B(net9),
    .Y(_04931_));
 sky130_fd_sc_hd__and3_1 _05803_ (.A(net55),
    .B(net9),
    .C(_04930_),
    .X(_04932_));
 sky130_fd_sc_hd__nand2b_1 _05804_ (.A_N(_04930_),
    .B(_04931_),
    .Y(_04933_));
 sky130_fd_sc_hd__xor2_1 _05805_ (.A(_04930_),
    .B(_04931_),
    .X(_04934_));
 sky130_fd_sc_hd__xnor2_1 _05806_ (.A(_04925_),
    .B(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__nand2_1 _05807_ (.A(net58),
    .B(net8),
    .Y(_04936_));
 sky130_fd_sc_hd__and3_1 _05808_ (.A(net58),
    .B(net8),
    .C(_04935_),
    .X(_04937_));
 sky130_fd_sc_hd__xnor2_1 _05809_ (.A(_04935_),
    .B(_04936_),
    .Y(_04938_));
 sky130_fd_sc_hd__xor2_1 _05810_ (.A(_04924_),
    .B(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__nand2_1 _05811_ (.A(net59),
    .B(net7),
    .Y(_04940_));
 sky130_fd_sc_hd__and3_1 _05812_ (.A(net59),
    .B(net7),
    .C(_04939_),
    .X(_04941_));
 sky130_fd_sc_hd__xnor2_1 _05813_ (.A(_04939_),
    .B(_04940_),
    .Y(_04942_));
 sky130_fd_sc_hd__xor2_1 _05814_ (.A(_04923_),
    .B(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__nand2_1 _05815_ (.A(net60),
    .B(net6),
    .Y(_04944_));
 sky130_fd_sc_hd__and3_1 _05816_ (.A(net60),
    .B(net6),
    .C(_04943_),
    .X(_04945_));
 sky130_fd_sc_hd__xnor2_1 _05817_ (.A(_04943_),
    .B(_04944_),
    .Y(_04946_));
 sky130_fd_sc_hd__xor2_1 _05818_ (.A(_04922_),
    .B(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__nand2_1 _05819_ (.A(net5),
    .B(net61),
    .Y(_04948_));
 sky130_fd_sc_hd__and3_1 _05820_ (.A(net5),
    .B(net61),
    .C(_04947_),
    .X(_04949_));
 sky130_fd_sc_hd__xnor2_1 _05821_ (.A(_04947_),
    .B(_04948_),
    .Y(_04950_));
 sky130_fd_sc_hd__xor2_1 _05822_ (.A(_04921_),
    .B(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__nand2_1 _05823_ (.A(net4),
    .B(net62),
    .Y(_04952_));
 sky130_fd_sc_hd__and3_1 _05824_ (.A(net4),
    .B(net62),
    .C(_04951_),
    .X(_04953_));
 sky130_fd_sc_hd__xnor2_1 _05825_ (.A(_04951_),
    .B(_04952_),
    .Y(_04954_));
 sky130_fd_sc_hd__xor2_1 _05826_ (.A(_04920_),
    .B(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__nand2_1 _05827_ (.A(net3),
    .B(net63),
    .Y(_04956_));
 sky130_fd_sc_hd__and3_1 _05828_ (.A(net3),
    .B(net63),
    .C(_04955_),
    .X(_04957_));
 sky130_fd_sc_hd__xnor2_1 _05829_ (.A(_04955_),
    .B(_04956_),
    .Y(_04958_));
 sky130_fd_sc_hd__xnor2_1 _05830_ (.A(_04919_),
    .B(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__nand2_1 _05831_ (.A(net64),
    .B(net2),
    .Y(_04960_));
 sky130_fd_sc_hd__nor2_1 _05832_ (.A(_04959_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__xor2_1 _05833_ (.A(_04959_),
    .B(_04960_),
    .X(_04962_));
 sky130_fd_sc_hd__xnor2_1 _05834_ (.A(_04918_),
    .B(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__nand2_1 _05835_ (.A(net34),
    .B(net32),
    .Y(_04964_));
 sky130_fd_sc_hd__nor2_1 _05836_ (.A(_04963_),
    .B(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hd__xor2_1 _05837_ (.A(_04963_),
    .B(_04964_),
    .X(_04966_));
 sky130_fd_sc_hd__xnor2_1 _05838_ (.A(_04917_),
    .B(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__nand2_1 _05839_ (.A(net35),
    .B(net31),
    .Y(_04968_));
 sky130_fd_sc_hd__nor2_1 _05840_ (.A(_04967_),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__xor2_1 _05841_ (.A(_04967_),
    .B(_04968_),
    .X(_04970_));
 sky130_fd_sc_hd__xnor2_1 _05842_ (.A(_04916_),
    .B(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__nand2_1 _05843_ (.A(net36),
    .B(net30),
    .Y(_04972_));
 sky130_fd_sc_hd__nor2_1 _05844_ (.A(_04971_),
    .B(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__xor2_1 _05845_ (.A(_04971_),
    .B(_04972_),
    .X(_04974_));
 sky130_fd_sc_hd__xnor2_1 _05846_ (.A(_04915_),
    .B(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hd__nand2_1 _05847_ (.A(net29),
    .B(net37),
    .Y(_04976_));
 sky130_fd_sc_hd__nor2_1 _05848_ (.A(_04975_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__xor2_1 _05849_ (.A(_04975_),
    .B(_04976_),
    .X(_04978_));
 sky130_fd_sc_hd__xnor2_1 _05850_ (.A(_04914_),
    .B(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__nand2_1 _05851_ (.A(net28),
    .B(net38),
    .Y(_04980_));
 sky130_fd_sc_hd__nor2_1 _05852_ (.A(_04979_),
    .B(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__xor2_1 _05853_ (.A(_04979_),
    .B(_04980_),
    .X(_04982_));
 sky130_fd_sc_hd__xnor2_1 _05854_ (.A(_04913_),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__nand2_1 _05855_ (.A(net27),
    .B(net39),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_1 _05856_ (.A(_04983_),
    .B(_00000_),
    .Y(_00001_));
 sky130_fd_sc_hd__xor2_1 _05857_ (.A(_04983_),
    .B(_00000_),
    .X(_00002_));
 sky130_fd_sc_hd__xnor2_1 _05858_ (.A(_04912_),
    .B(_00002_),
    .Y(_00003_));
 sky130_fd_sc_hd__nand2_1 _05859_ (.A(net26),
    .B(net40),
    .Y(_00004_));
 sky130_fd_sc_hd__nor2_1 _05860_ (.A(_00003_),
    .B(_00004_),
    .Y(_00005_));
 sky130_fd_sc_hd__xor2_1 _05861_ (.A(_00003_),
    .B(_00004_),
    .X(_00006_));
 sky130_fd_sc_hd__xnor2_1 _05862_ (.A(_04911_),
    .B(_00006_),
    .Y(_00007_));
 sky130_fd_sc_hd__nand2_1 _05863_ (.A(net23),
    .B(net41),
    .Y(_00008_));
 sky130_fd_sc_hd__nor2_1 _05864_ (.A(_00007_),
    .B(_00008_),
    .Y(_00009_));
 sky130_fd_sc_hd__xor2_1 _05865_ (.A(_00007_),
    .B(_00008_),
    .X(_00010_));
 sky130_fd_sc_hd__xnor2_1 _05866_ (.A(_04910_),
    .B(_00010_),
    .Y(_00011_));
 sky130_fd_sc_hd__nand2_1 _05867_ (.A(net12),
    .B(net42),
    .Y(_00012_));
 sky130_fd_sc_hd__nor2_1 _05868_ (.A(_00011_),
    .B(_00012_),
    .Y(_00013_));
 sky130_fd_sc_hd__xor2_1 _05869_ (.A(_00011_),
    .B(_00012_),
    .X(_00014_));
 sky130_fd_sc_hd__xor2_1 _05870_ (.A(_04908_),
    .B(_00014_),
    .X(_00015_));
 sky130_fd_sc_hd__and3_1 _05871_ (.A(net1),
    .B(net43),
    .C(_00015_),
    .X(_00016_));
 sky130_fd_sc_hd__a21oi_1 _05872_ (.A1(net1),
    .A2(net43),
    .B1(_00015_),
    .Y(_00017_));
 sky130_fd_sc_hd__nor2_1 _05873_ (.A(_00016_),
    .B(_00017_),
    .Y(\genblk2[18].rca.ripple_adders[19].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _05874_ (.A1(_04908_),
    .A2(_00014_),
    .B1(_00013_),
    .X(_00018_));
 sky130_fd_sc_hd__a21o_1 _05875_ (.A1(_04910_),
    .A2(_00010_),
    .B1(_00009_),
    .X(_00019_));
 sky130_fd_sc_hd__a21o_1 _05876_ (.A1(_04911_),
    .A2(_00006_),
    .B1(_00005_),
    .X(_00020_));
 sky130_fd_sc_hd__a21o_1 _05877_ (.A1(_04912_),
    .A2(_00002_),
    .B1(_00001_),
    .X(_00021_));
 sky130_fd_sc_hd__a21o_1 _05878_ (.A1(_04913_),
    .A2(_04982_),
    .B1(_04981_),
    .X(_00022_));
 sky130_fd_sc_hd__a21o_1 _05879_ (.A1(_04914_),
    .A2(_04978_),
    .B1(_04977_),
    .X(_00023_));
 sky130_fd_sc_hd__a21o_1 _05880_ (.A1(_04915_),
    .A2(_04974_),
    .B1(_04973_),
    .X(_00024_));
 sky130_fd_sc_hd__a21o_1 _05881_ (.A1(_04916_),
    .A2(_04970_),
    .B1(_04969_),
    .X(_00025_));
 sky130_fd_sc_hd__a21o_1 _05882_ (.A1(_04917_),
    .A2(_04966_),
    .B1(_04965_),
    .X(_00026_));
 sky130_fd_sc_hd__a21o_1 _05883_ (.A1(_04918_),
    .A2(_04962_),
    .B1(_04961_),
    .X(_00027_));
 sky130_fd_sc_hd__a21o_1 _05884_ (.A1(_04919_),
    .A2(_04958_),
    .B1(_04957_),
    .X(_00028_));
 sky130_fd_sc_hd__a21o_1 _05885_ (.A1(_04920_),
    .A2(_04954_),
    .B1(_04953_),
    .X(_00029_));
 sky130_fd_sc_hd__a21o_1 _05886_ (.A1(_04921_),
    .A2(_04950_),
    .B1(_04949_),
    .X(_00030_));
 sky130_fd_sc_hd__a21o_1 _05887_ (.A1(_04922_),
    .A2(_04946_),
    .B1(_04945_),
    .X(_00031_));
 sky130_fd_sc_hd__a21o_1 _05888_ (.A1(_04923_),
    .A2(_04942_),
    .B1(_04941_),
    .X(_00032_));
 sky130_fd_sc_hd__a21o_1 _05889_ (.A1(_04924_),
    .A2(_04938_),
    .B1(_04937_),
    .X(_00033_));
 sky130_fd_sc_hd__a21o_1 _05890_ (.A1(_04925_),
    .A2(_04933_),
    .B1(_04932_),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_1 _05891_ (.A1(net44),
    .A2(net11),
    .B1(net13),
    .B2(net33),
    .X(_00035_));
 sky130_fd_sc_hd__and3_1 _05892_ (.A(net44),
    .B(net11),
    .C(net13),
    .X(_00036_));
 sky130_fd_sc_hd__a21bo_1 _05893_ (.A1(net33),
    .A2(_00036_),
    .B1_N(_00035_),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_1 _05894_ (.A1(net33),
    .A2(_04927_),
    .B1(_04929_),
    .B2(_04926_),
    .X(_00038_));
 sky130_fd_sc_hd__xnor2_1 _05895_ (.A(_00037_),
    .B(_00038_),
    .Y(_00039_));
 sky130_fd_sc_hd__nand2_1 _05896_ (.A(net55),
    .B(net10),
    .Y(_00040_));
 sky130_fd_sc_hd__and3_1 _05897_ (.A(net55),
    .B(net10),
    .C(_00039_),
    .X(_00041_));
 sky130_fd_sc_hd__nand2b_1 _05898_ (.A_N(_00039_),
    .B(_00040_),
    .Y(_00042_));
 sky130_fd_sc_hd__xor2_1 _05899_ (.A(_00039_),
    .B(_00040_),
    .X(_00043_));
 sky130_fd_sc_hd__xnor2_1 _05900_ (.A(_00034_),
    .B(_00043_),
    .Y(_00044_));
 sky130_fd_sc_hd__nand2_1 _05901_ (.A(net58),
    .B(net9),
    .Y(_00045_));
 sky130_fd_sc_hd__and3_1 _05902_ (.A(net58),
    .B(net9),
    .C(_00044_),
    .X(_00046_));
 sky130_fd_sc_hd__xnor2_1 _05903_ (.A(_00044_),
    .B(_00045_),
    .Y(_00047_));
 sky130_fd_sc_hd__xor2_1 _05904_ (.A(_00033_),
    .B(_00047_),
    .X(_00048_));
 sky130_fd_sc_hd__nand2_1 _05905_ (.A(net59),
    .B(net8),
    .Y(_00049_));
 sky130_fd_sc_hd__and3_1 _05906_ (.A(net59),
    .B(net8),
    .C(_00048_),
    .X(_00050_));
 sky130_fd_sc_hd__xnor2_1 _05907_ (.A(_00048_),
    .B(_00049_),
    .Y(_00051_));
 sky130_fd_sc_hd__xor2_1 _05908_ (.A(_00032_),
    .B(_00051_),
    .X(_00052_));
 sky130_fd_sc_hd__nand2_1 _05909_ (.A(net60),
    .B(net7),
    .Y(_00053_));
 sky130_fd_sc_hd__and3_1 _05910_ (.A(net60),
    .B(net7),
    .C(_00052_),
    .X(_00054_));
 sky130_fd_sc_hd__xnor2_1 _05911_ (.A(_00052_),
    .B(_00053_),
    .Y(_00055_));
 sky130_fd_sc_hd__xor2_1 _05912_ (.A(_00031_),
    .B(_00055_),
    .X(_00056_));
 sky130_fd_sc_hd__nand2_1 _05913_ (.A(net61),
    .B(net6),
    .Y(_00057_));
 sky130_fd_sc_hd__and3_1 _05914_ (.A(net61),
    .B(net6),
    .C(_00056_),
    .X(_00058_));
 sky130_fd_sc_hd__xnor2_1 _05915_ (.A(_00056_),
    .B(_00057_),
    .Y(_00059_));
 sky130_fd_sc_hd__xor2_1 _05916_ (.A(_00030_),
    .B(_00059_),
    .X(_00060_));
 sky130_fd_sc_hd__nand2_1 _05917_ (.A(net5),
    .B(net62),
    .Y(_00061_));
 sky130_fd_sc_hd__and3_1 _05918_ (.A(net5),
    .B(net62),
    .C(_00060_),
    .X(_00062_));
 sky130_fd_sc_hd__xnor2_1 _05919_ (.A(_00060_),
    .B(_00061_),
    .Y(_00063_));
 sky130_fd_sc_hd__xor2_1 _05920_ (.A(_00029_),
    .B(_00063_),
    .X(_00064_));
 sky130_fd_sc_hd__nand2_1 _05921_ (.A(net4),
    .B(net63),
    .Y(_00065_));
 sky130_fd_sc_hd__and3_1 _05922_ (.A(net4),
    .B(net63),
    .C(_00064_),
    .X(_00066_));
 sky130_fd_sc_hd__xnor2_1 _05923_ (.A(_00064_),
    .B(_00065_),
    .Y(_00067_));
 sky130_fd_sc_hd__xnor2_1 _05924_ (.A(_00028_),
    .B(_00067_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand2_1 _05925_ (.A(net64),
    .B(net3),
    .Y(_00069_));
 sky130_fd_sc_hd__nor2_1 _05926_ (.A(_00068_),
    .B(_00069_),
    .Y(_00070_));
 sky130_fd_sc_hd__xor2_1 _05927_ (.A(_00068_),
    .B(_00069_),
    .X(_00071_));
 sky130_fd_sc_hd__xnor2_1 _05928_ (.A(_00027_),
    .B(_00071_),
    .Y(_00072_));
 sky130_fd_sc_hd__nand2_1 _05929_ (.A(net34),
    .B(net2),
    .Y(_00073_));
 sky130_fd_sc_hd__nor2_1 _05930_ (.A(_00072_),
    .B(_00073_),
    .Y(_00074_));
 sky130_fd_sc_hd__xor2_1 _05931_ (.A(_00072_),
    .B(_00073_),
    .X(_00075_));
 sky130_fd_sc_hd__xnor2_1 _05932_ (.A(_00026_),
    .B(_00075_),
    .Y(_00076_));
 sky130_fd_sc_hd__nand2_1 _05933_ (.A(net35),
    .B(net32),
    .Y(_00077_));
 sky130_fd_sc_hd__nor2_1 _05934_ (.A(_00076_),
    .B(_00077_),
    .Y(_00078_));
 sky130_fd_sc_hd__xor2_1 _05935_ (.A(_00076_),
    .B(_00077_),
    .X(_00079_));
 sky130_fd_sc_hd__xnor2_1 _05936_ (.A(_00025_),
    .B(_00079_),
    .Y(_00080_));
 sky130_fd_sc_hd__nand2_1 _05937_ (.A(net36),
    .B(net31),
    .Y(_00081_));
 sky130_fd_sc_hd__nor2_1 _05938_ (.A(_00080_),
    .B(_00081_),
    .Y(_00082_));
 sky130_fd_sc_hd__xor2_1 _05939_ (.A(_00080_),
    .B(_00081_),
    .X(_00083_));
 sky130_fd_sc_hd__xnor2_1 _05940_ (.A(_00024_),
    .B(_00083_),
    .Y(_00084_));
 sky130_fd_sc_hd__nand2_1 _05941_ (.A(net30),
    .B(net37),
    .Y(_00085_));
 sky130_fd_sc_hd__nor2_1 _05942_ (.A(_00084_),
    .B(_00085_),
    .Y(_00086_));
 sky130_fd_sc_hd__xor2_1 _05943_ (.A(_00084_),
    .B(_00085_),
    .X(_00087_));
 sky130_fd_sc_hd__xnor2_1 _05944_ (.A(_00023_),
    .B(_00087_),
    .Y(_00088_));
 sky130_fd_sc_hd__nand2_1 _05945_ (.A(net29),
    .B(net38),
    .Y(_00089_));
 sky130_fd_sc_hd__nor2_1 _05946_ (.A(_00088_),
    .B(_00089_),
    .Y(_00090_));
 sky130_fd_sc_hd__xor2_1 _05947_ (.A(_00088_),
    .B(_00089_),
    .X(_00091_));
 sky130_fd_sc_hd__xnor2_1 _05948_ (.A(_00022_),
    .B(_00091_),
    .Y(_00092_));
 sky130_fd_sc_hd__nand2_1 _05949_ (.A(net28),
    .B(net39),
    .Y(_00093_));
 sky130_fd_sc_hd__nor2_1 _05950_ (.A(_00092_),
    .B(_00093_),
    .Y(_00094_));
 sky130_fd_sc_hd__xor2_1 _05951_ (.A(_00092_),
    .B(_00093_),
    .X(_00095_));
 sky130_fd_sc_hd__xnor2_1 _05952_ (.A(_00021_),
    .B(_00095_),
    .Y(_00096_));
 sky130_fd_sc_hd__nand2_1 _05953_ (.A(net27),
    .B(net40),
    .Y(_00097_));
 sky130_fd_sc_hd__nor2_1 _05954_ (.A(_00096_),
    .B(_00097_),
    .Y(_00098_));
 sky130_fd_sc_hd__xor2_1 _05955_ (.A(_00096_),
    .B(_00097_),
    .X(_00099_));
 sky130_fd_sc_hd__xnor2_1 _05956_ (.A(_00020_),
    .B(_00099_),
    .Y(_00100_));
 sky130_fd_sc_hd__nand2_1 _05957_ (.A(net26),
    .B(net41),
    .Y(_00101_));
 sky130_fd_sc_hd__nor2_1 _05958_ (.A(_00100_),
    .B(_00101_),
    .Y(_00102_));
 sky130_fd_sc_hd__xor2_1 _05959_ (.A(_00100_),
    .B(_00101_),
    .X(_00103_));
 sky130_fd_sc_hd__xnor2_1 _05960_ (.A(_00019_),
    .B(_00103_),
    .Y(_00104_));
 sky130_fd_sc_hd__nand2_1 _05961_ (.A(net23),
    .B(net42),
    .Y(_00105_));
 sky130_fd_sc_hd__nor2_1 _05962_ (.A(_00104_),
    .B(_00105_),
    .Y(_00106_));
 sky130_fd_sc_hd__xor2_1 _05963_ (.A(_00104_),
    .B(_00105_),
    .X(_00107_));
 sky130_fd_sc_hd__xnor2_1 _05964_ (.A(_00018_),
    .B(_00107_),
    .Y(_00108_));
 sky130_fd_sc_hd__nand2_1 _05965_ (.A(net12),
    .B(net43),
    .Y(_00109_));
 sky130_fd_sc_hd__nor2_1 _05966_ (.A(_00108_),
    .B(_00109_),
    .Y(_00110_));
 sky130_fd_sc_hd__xor2_1 _05967_ (.A(_00108_),
    .B(_00109_),
    .X(_00111_));
 sky130_fd_sc_hd__xor2_1 _05968_ (.A(_00016_),
    .B(_00111_),
    .X(_00112_));
 sky130_fd_sc_hd__and3_1 _05969_ (.A(net1),
    .B(net45),
    .C(_00112_),
    .X(_00113_));
 sky130_fd_sc_hd__a21oi_1 _05970_ (.A1(net1),
    .A2(net45),
    .B1(_00112_),
    .Y(_00114_));
 sky130_fd_sc_hd__nor2_1 _05971_ (.A(_00113_),
    .B(_00114_),
    .Y(\genblk2[19].rca.ripple_adders[20].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _05972_ (.A1(_00016_),
    .A2(_00111_),
    .B1(_00110_),
    .X(_00115_));
 sky130_fd_sc_hd__a21o_1 _05973_ (.A1(_00018_),
    .A2(_00107_),
    .B1(_00106_),
    .X(_00116_));
 sky130_fd_sc_hd__a21o_1 _05974_ (.A1(_00019_),
    .A2(_00103_),
    .B1(_00102_),
    .X(_00117_));
 sky130_fd_sc_hd__a21o_1 _05975_ (.A1(_00020_),
    .A2(_00099_),
    .B1(_00098_),
    .X(_00118_));
 sky130_fd_sc_hd__a21o_1 _05976_ (.A1(_00021_),
    .A2(_00095_),
    .B1(_00094_),
    .X(_00119_));
 sky130_fd_sc_hd__a21o_1 _05977_ (.A1(_00022_),
    .A2(_00091_),
    .B1(_00090_),
    .X(_00120_));
 sky130_fd_sc_hd__a21o_1 _05978_ (.A1(_00023_),
    .A2(_00087_),
    .B1(_00086_),
    .X(_00121_));
 sky130_fd_sc_hd__a21o_1 _05979_ (.A1(_00024_),
    .A2(_00083_),
    .B1(_00082_),
    .X(_00122_));
 sky130_fd_sc_hd__a21o_1 _05980_ (.A1(_00025_),
    .A2(_00079_),
    .B1(_00078_),
    .X(_00123_));
 sky130_fd_sc_hd__a21o_1 _05981_ (.A1(_00026_),
    .A2(_00075_),
    .B1(_00074_),
    .X(_00124_));
 sky130_fd_sc_hd__a21o_1 _05982_ (.A1(_00027_),
    .A2(_00071_),
    .B1(_00070_),
    .X(_00125_));
 sky130_fd_sc_hd__a21o_1 _05983_ (.A1(_00028_),
    .A2(_00067_),
    .B1(_00066_),
    .X(_00126_));
 sky130_fd_sc_hd__a21o_1 _05984_ (.A1(_00029_),
    .A2(_00063_),
    .B1(_00062_),
    .X(_00127_));
 sky130_fd_sc_hd__a21o_1 _05985_ (.A1(_00030_),
    .A2(_00059_),
    .B1(_00058_),
    .X(_00128_));
 sky130_fd_sc_hd__a21o_1 _05986_ (.A1(_00031_),
    .A2(_00055_),
    .B1(_00054_),
    .X(_00129_));
 sky130_fd_sc_hd__a21o_1 _05987_ (.A1(_00032_),
    .A2(_00051_),
    .B1(_00050_),
    .X(_00130_));
 sky130_fd_sc_hd__a21o_1 _05988_ (.A1(_00033_),
    .A2(_00047_),
    .B1(_00046_),
    .X(_00131_));
 sky130_fd_sc_hd__a21o_1 _05989_ (.A1(_00034_),
    .A2(_00042_),
    .B1(_00041_),
    .X(_00132_));
 sky130_fd_sc_hd__a22o_1 _05990_ (.A1(net44),
    .A2(net13),
    .B1(net14),
    .B2(net33),
    .X(_00133_));
 sky130_fd_sc_hd__and3_1 _05991_ (.A(net44),
    .B(net13),
    .C(net14),
    .X(_00134_));
 sky130_fd_sc_hd__a21bo_1 _05992_ (.A1(net33),
    .A2(_00134_),
    .B1_N(_00133_),
    .X(_00135_));
 sky130_fd_sc_hd__a22o_1 _05993_ (.A1(net33),
    .A2(_00036_),
    .B1(_00038_),
    .B2(_00035_),
    .X(_00136_));
 sky130_fd_sc_hd__xnor2_1 _05994_ (.A(_00135_),
    .B(_00136_),
    .Y(_00137_));
 sky130_fd_sc_hd__nand2_1 _05995_ (.A(net55),
    .B(net11),
    .Y(_00138_));
 sky130_fd_sc_hd__and3_1 _05996_ (.A(net55),
    .B(net11),
    .C(_00137_),
    .X(_00139_));
 sky130_fd_sc_hd__nand2b_1 _05997_ (.A_N(_00137_),
    .B(_00138_),
    .Y(_00140_));
 sky130_fd_sc_hd__xor2_1 _05998_ (.A(_00137_),
    .B(_00138_),
    .X(_00141_));
 sky130_fd_sc_hd__xnor2_1 _05999_ (.A(_00132_),
    .B(_00141_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand2_1 _06000_ (.A(net58),
    .B(net10),
    .Y(_00143_));
 sky130_fd_sc_hd__and3_1 _06001_ (.A(net58),
    .B(net10),
    .C(_00142_),
    .X(_00144_));
 sky130_fd_sc_hd__xnor2_1 _06002_ (.A(_00142_),
    .B(_00143_),
    .Y(_00145_));
 sky130_fd_sc_hd__xor2_1 _06003_ (.A(_00131_),
    .B(_00145_),
    .X(_00146_));
 sky130_fd_sc_hd__nand2_1 _06004_ (.A(net59),
    .B(net9),
    .Y(_00147_));
 sky130_fd_sc_hd__and3_1 _06005_ (.A(net59),
    .B(net9),
    .C(_00146_),
    .X(_00148_));
 sky130_fd_sc_hd__xnor2_1 _06006_ (.A(_00146_),
    .B(_00147_),
    .Y(_00149_));
 sky130_fd_sc_hd__xor2_1 _06007_ (.A(_00130_),
    .B(_00149_),
    .X(_00150_));
 sky130_fd_sc_hd__nand2_1 _06008_ (.A(net60),
    .B(net8),
    .Y(_00151_));
 sky130_fd_sc_hd__and3_1 _06009_ (.A(net60),
    .B(net8),
    .C(_00150_),
    .X(_00152_));
 sky130_fd_sc_hd__xnor2_1 _06010_ (.A(_00150_),
    .B(_00151_),
    .Y(_00153_));
 sky130_fd_sc_hd__xor2_1 _06011_ (.A(_00129_),
    .B(_00153_),
    .X(_00154_));
 sky130_fd_sc_hd__nand2_1 _06012_ (.A(net61),
    .B(net7),
    .Y(_00155_));
 sky130_fd_sc_hd__and3_1 _06013_ (.A(net61),
    .B(net7),
    .C(_00154_),
    .X(_00156_));
 sky130_fd_sc_hd__xnor2_1 _06014_ (.A(_00154_),
    .B(_00155_),
    .Y(_00157_));
 sky130_fd_sc_hd__xor2_1 _06015_ (.A(_00128_),
    .B(_00157_),
    .X(_00158_));
 sky130_fd_sc_hd__nand2_1 _06016_ (.A(net62),
    .B(net6),
    .Y(_00159_));
 sky130_fd_sc_hd__and3_1 _06017_ (.A(net62),
    .B(net6),
    .C(_00158_),
    .X(_00160_));
 sky130_fd_sc_hd__xnor2_1 _06018_ (.A(_00158_),
    .B(_00159_),
    .Y(_00161_));
 sky130_fd_sc_hd__xor2_1 _06019_ (.A(_00127_),
    .B(_00161_),
    .X(_00162_));
 sky130_fd_sc_hd__nand2_1 _06020_ (.A(net5),
    .B(net63),
    .Y(_00163_));
 sky130_fd_sc_hd__and3_1 _06021_ (.A(net5),
    .B(net63),
    .C(_00162_),
    .X(_00164_));
 sky130_fd_sc_hd__xnor2_1 _06022_ (.A(_00162_),
    .B(_00163_),
    .Y(_00165_));
 sky130_fd_sc_hd__xnor2_1 _06023_ (.A(_00126_),
    .B(_00165_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand2_1 _06024_ (.A(net64),
    .B(net4),
    .Y(_00167_));
 sky130_fd_sc_hd__nor2_1 _06025_ (.A(_00166_),
    .B(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__xor2_1 _06026_ (.A(_00166_),
    .B(_00167_),
    .X(_00169_));
 sky130_fd_sc_hd__xnor2_1 _06027_ (.A(_00125_),
    .B(_00169_),
    .Y(_00170_));
 sky130_fd_sc_hd__nand2_1 _06028_ (.A(net34),
    .B(net3),
    .Y(_00171_));
 sky130_fd_sc_hd__nor2_1 _06029_ (.A(_00170_),
    .B(_00171_),
    .Y(_00172_));
 sky130_fd_sc_hd__xor2_1 _06030_ (.A(_00170_),
    .B(_00171_),
    .X(_00173_));
 sky130_fd_sc_hd__xnor2_1 _06031_ (.A(_00124_),
    .B(_00173_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _06032_ (.A(net35),
    .B(net2),
    .Y(_00175_));
 sky130_fd_sc_hd__nor2_1 _06033_ (.A(_00174_),
    .B(_00175_),
    .Y(_00176_));
 sky130_fd_sc_hd__xor2_1 _06034_ (.A(_00174_),
    .B(_00175_),
    .X(_00177_));
 sky130_fd_sc_hd__xnor2_1 _06035_ (.A(_00123_),
    .B(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _06036_ (.A(net36),
    .B(net32),
    .Y(_00179_));
 sky130_fd_sc_hd__nor2_1 _06037_ (.A(_00178_),
    .B(_00179_),
    .Y(_00180_));
 sky130_fd_sc_hd__xor2_1 _06038_ (.A(_00178_),
    .B(_00179_),
    .X(_00181_));
 sky130_fd_sc_hd__xnor2_1 _06039_ (.A(_00122_),
    .B(_00181_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand2_1 _06040_ (.A(net31),
    .B(net37),
    .Y(_00183_));
 sky130_fd_sc_hd__nor2_1 _06041_ (.A(_00182_),
    .B(_00183_),
    .Y(_00184_));
 sky130_fd_sc_hd__xor2_1 _06042_ (.A(_00182_),
    .B(_00183_),
    .X(_00185_));
 sky130_fd_sc_hd__xnor2_1 _06043_ (.A(_00121_),
    .B(_00185_),
    .Y(_00186_));
 sky130_fd_sc_hd__nand2_1 _06044_ (.A(net30),
    .B(net38),
    .Y(_00187_));
 sky130_fd_sc_hd__nor2_1 _06045_ (.A(_00186_),
    .B(_00187_),
    .Y(_00188_));
 sky130_fd_sc_hd__xor2_1 _06046_ (.A(_00186_),
    .B(_00187_),
    .X(_00189_));
 sky130_fd_sc_hd__xnor2_1 _06047_ (.A(_00120_),
    .B(_00189_),
    .Y(_00190_));
 sky130_fd_sc_hd__nand2_1 _06048_ (.A(net29),
    .B(net39),
    .Y(_00191_));
 sky130_fd_sc_hd__nor2_1 _06049_ (.A(_00190_),
    .B(_00191_),
    .Y(_00192_));
 sky130_fd_sc_hd__xor2_1 _06050_ (.A(_00190_),
    .B(_00191_),
    .X(_00193_));
 sky130_fd_sc_hd__xnor2_1 _06051_ (.A(_00119_),
    .B(_00193_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _06052_ (.A(net28),
    .B(net40),
    .Y(_00195_));
 sky130_fd_sc_hd__nor2_1 _06053_ (.A(_00194_),
    .B(_00195_),
    .Y(_00196_));
 sky130_fd_sc_hd__xor2_1 _06054_ (.A(_00194_),
    .B(_00195_),
    .X(_00197_));
 sky130_fd_sc_hd__xnor2_1 _06055_ (.A(_00118_),
    .B(_00197_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _06056_ (.A(net27),
    .B(net41),
    .Y(_00199_));
 sky130_fd_sc_hd__nor2_1 _06057_ (.A(_00198_),
    .B(_00199_),
    .Y(_00200_));
 sky130_fd_sc_hd__xor2_1 _06058_ (.A(_00198_),
    .B(_00199_),
    .X(_00201_));
 sky130_fd_sc_hd__xnor2_1 _06059_ (.A(_00117_),
    .B(_00201_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand2_1 _06060_ (.A(net26),
    .B(net42),
    .Y(_00203_));
 sky130_fd_sc_hd__nor2_1 _06061_ (.A(_00202_),
    .B(_00203_),
    .Y(_00204_));
 sky130_fd_sc_hd__xor2_1 _06062_ (.A(_00202_),
    .B(_00203_),
    .X(_00205_));
 sky130_fd_sc_hd__xnor2_1 _06063_ (.A(_00116_),
    .B(_00205_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _06064_ (.A(net23),
    .B(net43),
    .Y(_00207_));
 sky130_fd_sc_hd__nor2_1 _06065_ (.A(_00206_),
    .B(_00207_),
    .Y(_00208_));
 sky130_fd_sc_hd__xor2_1 _06066_ (.A(_00206_),
    .B(_00207_),
    .X(_00209_));
 sky130_fd_sc_hd__xnor2_1 _06067_ (.A(_00115_),
    .B(_00209_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _06068_ (.A(net12),
    .B(net45),
    .Y(_00211_));
 sky130_fd_sc_hd__nor2_1 _06069_ (.A(_00210_),
    .B(_00211_),
    .Y(_00212_));
 sky130_fd_sc_hd__xor2_1 _06070_ (.A(_00210_),
    .B(_00211_),
    .X(_00213_));
 sky130_fd_sc_hd__xor2_1 _06071_ (.A(_00113_),
    .B(_00213_),
    .X(_00214_));
 sky130_fd_sc_hd__and3_1 _06072_ (.A(net1),
    .B(net46),
    .C(_00214_),
    .X(_00215_));
 sky130_fd_sc_hd__a21oi_1 _06073_ (.A1(net1),
    .A2(net46),
    .B1(_00214_),
    .Y(_00216_));
 sky130_fd_sc_hd__nor2_1 _06074_ (.A(_00215_),
    .B(_00216_),
    .Y(\genblk2[20].rca.ripple_adders[21].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _06075_ (.A1(_00113_),
    .A2(_00213_),
    .B1(_00212_),
    .X(_00217_));
 sky130_fd_sc_hd__a21o_1 _06076_ (.A1(_00115_),
    .A2(_00209_),
    .B1(_00208_),
    .X(_00218_));
 sky130_fd_sc_hd__a21o_1 _06077_ (.A1(_00116_),
    .A2(_00205_),
    .B1(_00204_),
    .X(_00219_));
 sky130_fd_sc_hd__a21o_1 _06078_ (.A1(_00117_),
    .A2(_00201_),
    .B1(_00200_),
    .X(_00220_));
 sky130_fd_sc_hd__a21o_1 _06079_ (.A1(_00118_),
    .A2(_00197_),
    .B1(_00196_),
    .X(_00221_));
 sky130_fd_sc_hd__a21o_1 _06080_ (.A1(_00119_),
    .A2(_00193_),
    .B1(_00192_),
    .X(_00222_));
 sky130_fd_sc_hd__a21o_1 _06081_ (.A1(_00120_),
    .A2(_00189_),
    .B1(_00188_),
    .X(_00223_));
 sky130_fd_sc_hd__a21o_1 _06082_ (.A1(_00121_),
    .A2(_00185_),
    .B1(_00184_),
    .X(_00224_));
 sky130_fd_sc_hd__a21o_1 _06083_ (.A1(_00122_),
    .A2(_00181_),
    .B1(_00180_),
    .X(_00225_));
 sky130_fd_sc_hd__a21o_1 _06084_ (.A1(_00123_),
    .A2(_00177_),
    .B1(_00176_),
    .X(_00226_));
 sky130_fd_sc_hd__a21o_1 _06085_ (.A1(_00124_),
    .A2(_00173_),
    .B1(_00172_),
    .X(_00227_));
 sky130_fd_sc_hd__a21o_1 _06086_ (.A1(_00125_),
    .A2(_00169_),
    .B1(_00168_),
    .X(_00228_));
 sky130_fd_sc_hd__a21o_1 _06087_ (.A1(_00126_),
    .A2(_00165_),
    .B1(_00164_),
    .X(_00229_));
 sky130_fd_sc_hd__a21o_1 _06088_ (.A1(_00127_),
    .A2(_00161_),
    .B1(_00160_),
    .X(_00230_));
 sky130_fd_sc_hd__a21o_1 _06089_ (.A1(_00128_),
    .A2(_00157_),
    .B1(_00156_),
    .X(_00231_));
 sky130_fd_sc_hd__a21o_1 _06090_ (.A1(_00129_),
    .A2(_00153_),
    .B1(_00152_),
    .X(_00232_));
 sky130_fd_sc_hd__a21o_1 _06091_ (.A1(_00130_),
    .A2(_00149_),
    .B1(_00148_),
    .X(_00233_));
 sky130_fd_sc_hd__a21o_1 _06092_ (.A1(_00131_),
    .A2(_00145_),
    .B1(_00144_),
    .X(_00234_));
 sky130_fd_sc_hd__a21o_1 _06093_ (.A1(_00132_),
    .A2(_00140_),
    .B1(_00139_),
    .X(_00235_));
 sky130_fd_sc_hd__a22o_1 _06094_ (.A1(net44),
    .A2(net14),
    .B1(net15),
    .B2(net33),
    .X(_00236_));
 sky130_fd_sc_hd__and3_1 _06095_ (.A(net44),
    .B(net14),
    .C(net15),
    .X(_00237_));
 sky130_fd_sc_hd__a21bo_1 _06096_ (.A1(net33),
    .A2(_00237_),
    .B1_N(_00236_),
    .X(_00238_));
 sky130_fd_sc_hd__a22o_1 _06097_ (.A1(net33),
    .A2(_00134_),
    .B1(_00136_),
    .B2(_00133_),
    .X(_00239_));
 sky130_fd_sc_hd__xnor2_1 _06098_ (.A(_00238_),
    .B(_00239_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _06099_ (.A(net55),
    .B(net13),
    .Y(_00241_));
 sky130_fd_sc_hd__and3_1 _06100_ (.A(net55),
    .B(net13),
    .C(_00240_),
    .X(_00242_));
 sky130_fd_sc_hd__nand2b_1 _06101_ (.A_N(_00240_),
    .B(_00241_),
    .Y(_00243_));
 sky130_fd_sc_hd__xor2_1 _06102_ (.A(_00240_),
    .B(_00241_),
    .X(_00244_));
 sky130_fd_sc_hd__xnor2_1 _06103_ (.A(_00235_),
    .B(_00244_),
    .Y(_00245_));
 sky130_fd_sc_hd__nand2_1 _06104_ (.A(net58),
    .B(net11),
    .Y(_00246_));
 sky130_fd_sc_hd__and3_1 _06105_ (.A(net58),
    .B(net11),
    .C(_00245_),
    .X(_00247_));
 sky130_fd_sc_hd__xnor2_1 _06106_ (.A(_00245_),
    .B(_00246_),
    .Y(_00248_));
 sky130_fd_sc_hd__xor2_1 _06107_ (.A(_00234_),
    .B(_00248_),
    .X(_00249_));
 sky130_fd_sc_hd__nand2_1 _06108_ (.A(net59),
    .B(net10),
    .Y(_00250_));
 sky130_fd_sc_hd__and3_1 _06109_ (.A(net59),
    .B(net10),
    .C(_00249_),
    .X(_00251_));
 sky130_fd_sc_hd__xnor2_1 _06110_ (.A(_00249_),
    .B(_00250_),
    .Y(_00252_));
 sky130_fd_sc_hd__xor2_1 _06111_ (.A(_00233_),
    .B(_00252_),
    .X(_00253_));
 sky130_fd_sc_hd__nand2_1 _06112_ (.A(net60),
    .B(net9),
    .Y(_00254_));
 sky130_fd_sc_hd__and3_1 _06113_ (.A(net60),
    .B(net9),
    .C(_00253_),
    .X(_00255_));
 sky130_fd_sc_hd__xnor2_1 _06114_ (.A(_00253_),
    .B(_00254_),
    .Y(_00256_));
 sky130_fd_sc_hd__xor2_1 _06115_ (.A(_00232_),
    .B(_00256_),
    .X(_00257_));
 sky130_fd_sc_hd__nand2_1 _06116_ (.A(net61),
    .B(net8),
    .Y(_00258_));
 sky130_fd_sc_hd__and3_1 _06117_ (.A(net61),
    .B(net8),
    .C(_00257_),
    .X(_00259_));
 sky130_fd_sc_hd__xnor2_1 _06118_ (.A(_00257_),
    .B(_00258_),
    .Y(_00260_));
 sky130_fd_sc_hd__xor2_1 _06119_ (.A(_00231_),
    .B(_00260_),
    .X(_00261_));
 sky130_fd_sc_hd__nand2_1 _06120_ (.A(net62),
    .B(net7),
    .Y(_00262_));
 sky130_fd_sc_hd__and3_1 _06121_ (.A(net62),
    .B(net7),
    .C(_00261_),
    .X(_00263_));
 sky130_fd_sc_hd__xnor2_1 _06122_ (.A(_00261_),
    .B(_00262_),
    .Y(_00264_));
 sky130_fd_sc_hd__xnor2_1 _06123_ (.A(_00230_),
    .B(_00264_),
    .Y(_00265_));
 sky130_fd_sc_hd__nand2_1 _06124_ (.A(net63),
    .B(net6),
    .Y(_00266_));
 sky130_fd_sc_hd__nor2_1 _06125_ (.A(_00265_),
    .B(_00266_),
    .Y(_00267_));
 sky130_fd_sc_hd__xor2_1 _06126_ (.A(_00265_),
    .B(_00266_),
    .X(_00268_));
 sky130_fd_sc_hd__xnor2_1 _06127_ (.A(_00229_),
    .B(_00268_),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_1 _06128_ (.A(net64),
    .B(net5),
    .Y(_00270_));
 sky130_fd_sc_hd__nor2_1 _06129_ (.A(_00269_),
    .B(_00270_),
    .Y(_00271_));
 sky130_fd_sc_hd__xor2_1 _06130_ (.A(_00269_),
    .B(_00270_),
    .X(_00272_));
 sky130_fd_sc_hd__xnor2_1 _06131_ (.A(_00228_),
    .B(_00272_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _06132_ (.A(net34),
    .B(net4),
    .Y(_00274_));
 sky130_fd_sc_hd__nor2_1 _06133_ (.A(_00273_),
    .B(_00274_),
    .Y(_00275_));
 sky130_fd_sc_hd__xor2_1 _06134_ (.A(_00273_),
    .B(_00274_),
    .X(_00276_));
 sky130_fd_sc_hd__xnor2_1 _06135_ (.A(_00227_),
    .B(_00276_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _06136_ (.A(net35),
    .B(net3),
    .Y(_00278_));
 sky130_fd_sc_hd__nor2_1 _06137_ (.A(_00277_),
    .B(_00278_),
    .Y(_00279_));
 sky130_fd_sc_hd__xor2_1 _06138_ (.A(_00277_),
    .B(_00278_),
    .X(_00280_));
 sky130_fd_sc_hd__xnor2_1 _06139_ (.A(_00226_),
    .B(_00280_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_1 _06140_ (.A(net36),
    .B(net2),
    .Y(_00282_));
 sky130_fd_sc_hd__nor2_1 _06141_ (.A(_00281_),
    .B(_00282_),
    .Y(_00283_));
 sky130_fd_sc_hd__xor2_1 _06142_ (.A(_00281_),
    .B(_00282_),
    .X(_00284_));
 sky130_fd_sc_hd__xnor2_1 _06143_ (.A(_00225_),
    .B(_00284_),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _06144_ (.A(net32),
    .B(net37),
    .Y(_00286_));
 sky130_fd_sc_hd__nor2_1 _06145_ (.A(_00285_),
    .B(_00286_),
    .Y(_00288_));
 sky130_fd_sc_hd__xor2_1 _06146_ (.A(_00285_),
    .B(_00286_),
    .X(_00289_));
 sky130_fd_sc_hd__xnor2_1 _06147_ (.A(_00224_),
    .B(_00289_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _06148_ (.A(net31),
    .B(net38),
    .Y(_00291_));
 sky130_fd_sc_hd__nor2_1 _06149_ (.A(_00290_),
    .B(_00291_),
    .Y(_00292_));
 sky130_fd_sc_hd__xor2_1 _06150_ (.A(_00290_),
    .B(_00291_),
    .X(_00293_));
 sky130_fd_sc_hd__xnor2_1 _06151_ (.A(_00223_),
    .B(_00293_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _06152_ (.A(net30),
    .B(net39),
    .Y(_00295_));
 sky130_fd_sc_hd__nor2_1 _06153_ (.A(_00294_),
    .B(_00295_),
    .Y(_00296_));
 sky130_fd_sc_hd__xor2_1 _06154_ (.A(_00294_),
    .B(_00295_),
    .X(_00297_));
 sky130_fd_sc_hd__xnor2_1 _06155_ (.A(_00222_),
    .B(_00297_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand2_1 _06156_ (.A(net29),
    .B(net40),
    .Y(_00300_));
 sky130_fd_sc_hd__nor2_1 _06157_ (.A(_00299_),
    .B(_00300_),
    .Y(_00301_));
 sky130_fd_sc_hd__xor2_1 _06158_ (.A(_00299_),
    .B(_00300_),
    .X(_00302_));
 sky130_fd_sc_hd__xnor2_1 _06159_ (.A(_00221_),
    .B(_00302_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _06160_ (.A(net28),
    .B(net41),
    .Y(_00304_));
 sky130_fd_sc_hd__nor2_1 _06161_ (.A(_00303_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__xor2_1 _06162_ (.A(_00303_),
    .B(_00304_),
    .X(_00306_));
 sky130_fd_sc_hd__xnor2_1 _06163_ (.A(_00220_),
    .B(_00306_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_1 _06164_ (.A(net27),
    .B(net42),
    .Y(_00308_));
 sky130_fd_sc_hd__nor2_1 _06165_ (.A(_00307_),
    .B(_00308_),
    .Y(_00310_));
 sky130_fd_sc_hd__xor2_1 _06166_ (.A(_00307_),
    .B(_00308_),
    .X(_00311_));
 sky130_fd_sc_hd__xnor2_1 _06167_ (.A(_00219_),
    .B(_00311_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _06168_ (.A(net26),
    .B(net43),
    .Y(_00313_));
 sky130_fd_sc_hd__nor2_1 _06169_ (.A(_00312_),
    .B(_00313_),
    .Y(_00314_));
 sky130_fd_sc_hd__xor2_1 _06170_ (.A(_00312_),
    .B(_00313_),
    .X(_00315_));
 sky130_fd_sc_hd__xnor2_1 _06171_ (.A(_00218_),
    .B(_00315_),
    .Y(_00316_));
 sky130_fd_sc_hd__nand2_1 _06172_ (.A(net23),
    .B(net45),
    .Y(_00317_));
 sky130_fd_sc_hd__nor2_1 _06173_ (.A(_00316_),
    .B(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__xor2_1 _06174_ (.A(_00316_),
    .B(_00317_),
    .X(_00319_));
 sky130_fd_sc_hd__xnor2_1 _06175_ (.A(_00217_),
    .B(_00319_),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _06176_ (.A(net12),
    .B(net46),
    .Y(_00321_));
 sky130_fd_sc_hd__nor2_1 _06177_ (.A(_00320_),
    .B(_00321_),
    .Y(_00322_));
 sky130_fd_sc_hd__xor2_1 _06178_ (.A(_00320_),
    .B(_00321_),
    .X(_00323_));
 sky130_fd_sc_hd__xor2_1 _06179_ (.A(_00215_),
    .B(_00323_),
    .X(_00324_));
 sky130_fd_sc_hd__and3_1 _06180_ (.A(net1),
    .B(net47),
    .C(_00324_),
    .X(_00325_));
 sky130_fd_sc_hd__a21oi_1 _06181_ (.A1(net1),
    .A2(net47),
    .B1(_00324_),
    .Y(_00326_));
 sky130_fd_sc_hd__nor2_1 _06182_ (.A(_00325_),
    .B(_00326_),
    .Y(\genblk2[21].rca.ripple_adders[22].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _06183_ (.A1(_00215_),
    .A2(_00323_),
    .B1(_00322_),
    .X(_00327_));
 sky130_fd_sc_hd__a21o_1 _06184_ (.A1(_00217_),
    .A2(_00319_),
    .B1(_00318_),
    .X(_00328_));
 sky130_fd_sc_hd__a21o_1 _06185_ (.A1(_00218_),
    .A2(_00315_),
    .B1(_00314_),
    .X(_00330_));
 sky130_fd_sc_hd__a21o_1 _06186_ (.A1(_00219_),
    .A2(_00311_),
    .B1(_00310_),
    .X(_00331_));
 sky130_fd_sc_hd__a21o_1 _06187_ (.A1(_00220_),
    .A2(_00306_),
    .B1(_00305_),
    .X(_00332_));
 sky130_fd_sc_hd__a21o_1 _06188_ (.A1(_00221_),
    .A2(_00302_),
    .B1(_00301_),
    .X(_00333_));
 sky130_fd_sc_hd__a21o_1 _06189_ (.A1(_00222_),
    .A2(_00297_),
    .B1(_00296_),
    .X(_00334_));
 sky130_fd_sc_hd__a21o_1 _06190_ (.A1(_00223_),
    .A2(_00293_),
    .B1(_00292_),
    .X(_00335_));
 sky130_fd_sc_hd__a21o_1 _06191_ (.A1(_00224_),
    .A2(_00289_),
    .B1(_00288_),
    .X(_00336_));
 sky130_fd_sc_hd__a21o_1 _06192_ (.A1(_00225_),
    .A2(_00284_),
    .B1(_00283_),
    .X(_00337_));
 sky130_fd_sc_hd__a21o_1 _06193_ (.A1(_00226_),
    .A2(_00280_),
    .B1(_00279_),
    .X(_00338_));
 sky130_fd_sc_hd__a21o_1 _06194_ (.A1(_00227_),
    .A2(_00276_),
    .B1(_00275_),
    .X(_00339_));
 sky130_fd_sc_hd__a21o_1 _06195_ (.A1(_00228_),
    .A2(_00272_),
    .B1(_00271_),
    .X(_00341_));
 sky130_fd_sc_hd__a21o_1 _06196_ (.A1(_00229_),
    .A2(_00268_),
    .B1(_00267_),
    .X(_00342_));
 sky130_fd_sc_hd__a21o_1 _06197_ (.A1(_00230_),
    .A2(_00264_),
    .B1(_00263_),
    .X(_00343_));
 sky130_fd_sc_hd__a21o_1 _06198_ (.A1(_00231_),
    .A2(_00260_),
    .B1(_00259_),
    .X(_00344_));
 sky130_fd_sc_hd__a21o_1 _06199_ (.A1(_00232_),
    .A2(_00256_),
    .B1(_00255_),
    .X(_00345_));
 sky130_fd_sc_hd__a21o_1 _06200_ (.A1(_00233_),
    .A2(_00252_),
    .B1(_00251_),
    .X(_00346_));
 sky130_fd_sc_hd__a21o_1 _06201_ (.A1(_00234_),
    .A2(_00248_),
    .B1(_00247_),
    .X(_00347_));
 sky130_fd_sc_hd__a21o_1 _06202_ (.A1(_00235_),
    .A2(_00243_),
    .B1(_00242_),
    .X(_00348_));
 sky130_fd_sc_hd__a22o_1 _06203_ (.A1(net44),
    .A2(net15),
    .B1(net16),
    .B2(net33),
    .X(_00349_));
 sky130_fd_sc_hd__and3_1 _06204_ (.A(net44),
    .B(net15),
    .C(net16),
    .X(_00350_));
 sky130_fd_sc_hd__a21bo_1 _06205_ (.A1(net33),
    .A2(_00350_),
    .B1_N(_00349_),
    .X(_00352_));
 sky130_fd_sc_hd__a22o_1 _06206_ (.A1(net33),
    .A2(_00237_),
    .B1(_00239_),
    .B2(_00236_),
    .X(_00353_));
 sky130_fd_sc_hd__xnor2_1 _06207_ (.A(_00352_),
    .B(_00353_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2_1 _06208_ (.A(net55),
    .B(net14),
    .Y(_00355_));
 sky130_fd_sc_hd__and3_1 _06209_ (.A(net55),
    .B(net14),
    .C(_00354_),
    .X(_00356_));
 sky130_fd_sc_hd__nand2b_1 _06210_ (.A_N(_00354_),
    .B(_00355_),
    .Y(_00357_));
 sky130_fd_sc_hd__xor2_1 _06211_ (.A(_00354_),
    .B(_00355_),
    .X(_00358_));
 sky130_fd_sc_hd__xnor2_1 _06212_ (.A(_00348_),
    .B(_00358_),
    .Y(_00359_));
 sky130_fd_sc_hd__nand2_1 _06213_ (.A(net58),
    .B(net13),
    .Y(_00360_));
 sky130_fd_sc_hd__and3_1 _06214_ (.A(net58),
    .B(net13),
    .C(_00359_),
    .X(_00361_));
 sky130_fd_sc_hd__xnor2_1 _06215_ (.A(_00359_),
    .B(_00360_),
    .Y(_00363_));
 sky130_fd_sc_hd__xor2_1 _06216_ (.A(_00347_),
    .B(_00363_),
    .X(_00364_));
 sky130_fd_sc_hd__nand2_1 _06217_ (.A(net59),
    .B(net11),
    .Y(_00365_));
 sky130_fd_sc_hd__and3_1 _06218_ (.A(net59),
    .B(net11),
    .C(_00364_),
    .X(_00366_));
 sky130_fd_sc_hd__xnor2_1 _06219_ (.A(_00364_),
    .B(_00365_),
    .Y(_00367_));
 sky130_fd_sc_hd__xor2_1 _06220_ (.A(_00346_),
    .B(_00367_),
    .X(_00368_));
 sky130_fd_sc_hd__nand2_1 _06221_ (.A(net60),
    .B(net10),
    .Y(_00369_));
 sky130_fd_sc_hd__and3_1 _06222_ (.A(net60),
    .B(net10),
    .C(_00368_),
    .X(_00370_));
 sky130_fd_sc_hd__xnor2_1 _06223_ (.A(_00368_),
    .B(_00369_),
    .Y(_00371_));
 sky130_fd_sc_hd__xor2_1 _06224_ (.A(_00345_),
    .B(_00371_),
    .X(_00372_));
 sky130_fd_sc_hd__nand2_1 _06225_ (.A(net61),
    .B(net9),
    .Y(_00374_));
 sky130_fd_sc_hd__and3_1 _06226_ (.A(net61),
    .B(net9),
    .C(_00372_),
    .X(_00375_));
 sky130_fd_sc_hd__xnor2_1 _06227_ (.A(_00372_),
    .B(_00374_),
    .Y(_00376_));
 sky130_fd_sc_hd__xor2_1 _06228_ (.A(_00344_),
    .B(_00376_),
    .X(_00377_));
 sky130_fd_sc_hd__nand2_1 _06229_ (.A(net62),
    .B(net8),
    .Y(_00378_));
 sky130_fd_sc_hd__and3_1 _06230_ (.A(net62),
    .B(net8),
    .C(_00377_),
    .X(_00379_));
 sky130_fd_sc_hd__xnor2_1 _06231_ (.A(_00377_),
    .B(_00378_),
    .Y(_00380_));
 sky130_fd_sc_hd__xnor2_1 _06232_ (.A(_00343_),
    .B(_00380_),
    .Y(_00381_));
 sky130_fd_sc_hd__nand2_1 _06233_ (.A(net63),
    .B(net7),
    .Y(_00382_));
 sky130_fd_sc_hd__nor2_1 _06234_ (.A(_00381_),
    .B(_00382_),
    .Y(_00383_));
 sky130_fd_sc_hd__xor2_1 _06235_ (.A(_00381_),
    .B(_00382_),
    .X(_00385_));
 sky130_fd_sc_hd__xnor2_1 _06236_ (.A(_00342_),
    .B(_00385_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _06237_ (.A(net64),
    .B(net6),
    .Y(_00387_));
 sky130_fd_sc_hd__nor2_1 _06238_ (.A(_00386_),
    .B(_00387_),
    .Y(_00388_));
 sky130_fd_sc_hd__xor2_1 _06239_ (.A(_00386_),
    .B(_00387_),
    .X(_00389_));
 sky130_fd_sc_hd__xnor2_1 _06240_ (.A(_00341_),
    .B(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _06241_ (.A(net34),
    .B(net5),
    .Y(_00391_));
 sky130_fd_sc_hd__nor2_1 _06242_ (.A(_00390_),
    .B(_00391_),
    .Y(_00392_));
 sky130_fd_sc_hd__xor2_1 _06243_ (.A(_00390_),
    .B(_00391_),
    .X(_00393_));
 sky130_fd_sc_hd__xnor2_1 _06244_ (.A(_00339_),
    .B(_00393_),
    .Y(_00394_));
 sky130_fd_sc_hd__nand2_1 _06245_ (.A(net35),
    .B(net4),
    .Y(_00396_));
 sky130_fd_sc_hd__nor2_1 _06246_ (.A(_00394_),
    .B(_00396_),
    .Y(_00397_));
 sky130_fd_sc_hd__xor2_1 _06247_ (.A(_00394_),
    .B(_00396_),
    .X(_00398_));
 sky130_fd_sc_hd__xnor2_1 _06248_ (.A(_00338_),
    .B(_00398_),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _06249_ (.A(net36),
    .B(net3),
    .Y(_00400_));
 sky130_fd_sc_hd__nor2_1 _06250_ (.A(_00399_),
    .B(_00400_),
    .Y(_00401_));
 sky130_fd_sc_hd__xor2_1 _06251_ (.A(_00399_),
    .B(_00400_),
    .X(_00402_));
 sky130_fd_sc_hd__xnor2_1 _06252_ (.A(_00337_),
    .B(_00402_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _06253_ (.A(net2),
    .B(net37),
    .Y(_00404_));
 sky130_fd_sc_hd__nor2_1 _06254_ (.A(_00403_),
    .B(_00404_),
    .Y(_00405_));
 sky130_fd_sc_hd__xor2_1 _06255_ (.A(_00403_),
    .B(_00404_),
    .X(_00407_));
 sky130_fd_sc_hd__xnor2_1 _06256_ (.A(_00336_),
    .B(_00407_),
    .Y(_00408_));
 sky130_fd_sc_hd__nand2_1 _06257_ (.A(net32),
    .B(net38),
    .Y(_00409_));
 sky130_fd_sc_hd__nor2_1 _06258_ (.A(_00408_),
    .B(_00409_),
    .Y(_00410_));
 sky130_fd_sc_hd__xor2_1 _06259_ (.A(_00408_),
    .B(_00409_),
    .X(_00411_));
 sky130_fd_sc_hd__xnor2_1 _06260_ (.A(_00335_),
    .B(_00411_),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_1 _06261_ (.A(net31),
    .B(net39),
    .Y(_00413_));
 sky130_fd_sc_hd__nor2_1 _06262_ (.A(_00412_),
    .B(_00413_),
    .Y(_00414_));
 sky130_fd_sc_hd__xor2_1 _06263_ (.A(_00412_),
    .B(_00413_),
    .X(_00415_));
 sky130_fd_sc_hd__xnor2_1 _06264_ (.A(_00334_),
    .B(_00415_),
    .Y(_00416_));
 sky130_fd_sc_hd__nand2_1 _06265_ (.A(net30),
    .B(net40),
    .Y(_00418_));
 sky130_fd_sc_hd__nor2_1 _06266_ (.A(_00416_),
    .B(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__xor2_1 _06267_ (.A(_00416_),
    .B(_00418_),
    .X(_00420_));
 sky130_fd_sc_hd__xnor2_1 _06268_ (.A(_00333_),
    .B(_00420_),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _06269_ (.A(net29),
    .B(net41),
    .Y(_00422_));
 sky130_fd_sc_hd__nor2_1 _06270_ (.A(_00421_),
    .B(_00422_),
    .Y(_00423_));
 sky130_fd_sc_hd__xor2_1 _06271_ (.A(_00421_),
    .B(_00422_),
    .X(_00424_));
 sky130_fd_sc_hd__xnor2_1 _06272_ (.A(_00332_),
    .B(_00424_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _06273_ (.A(net28),
    .B(net42),
    .Y(_00426_));
 sky130_fd_sc_hd__nor2_1 _06274_ (.A(_00425_),
    .B(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__xor2_1 _06275_ (.A(_00425_),
    .B(_00426_),
    .X(_00429_));
 sky130_fd_sc_hd__xnor2_1 _06276_ (.A(_00331_),
    .B(_00429_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _06277_ (.A(net27),
    .B(net43),
    .Y(_00431_));
 sky130_fd_sc_hd__nor2_1 _06278_ (.A(_00430_),
    .B(_00431_),
    .Y(_00432_));
 sky130_fd_sc_hd__xor2_1 _06279_ (.A(_00430_),
    .B(_00431_),
    .X(_00433_));
 sky130_fd_sc_hd__xnor2_1 _06280_ (.A(_00330_),
    .B(_00433_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _06281_ (.A(net26),
    .B(net45),
    .Y(_00435_));
 sky130_fd_sc_hd__nor2_1 _06282_ (.A(_00434_),
    .B(_00435_),
    .Y(_00436_));
 sky130_fd_sc_hd__xor2_1 _06283_ (.A(_00434_),
    .B(_00435_),
    .X(_00437_));
 sky130_fd_sc_hd__xnor2_1 _06284_ (.A(_00328_),
    .B(_00437_),
    .Y(_00438_));
 sky130_fd_sc_hd__nand2_1 _06285_ (.A(net23),
    .B(net46),
    .Y(_00440_));
 sky130_fd_sc_hd__nor2_1 _06286_ (.A(_00438_),
    .B(_00440_),
    .Y(_00441_));
 sky130_fd_sc_hd__xor2_1 _06287_ (.A(_00438_),
    .B(_00440_),
    .X(_00442_));
 sky130_fd_sc_hd__xnor2_1 _06288_ (.A(_00327_),
    .B(_00442_),
    .Y(_00443_));
 sky130_fd_sc_hd__nand2_1 _06289_ (.A(net12),
    .B(net47),
    .Y(_00444_));
 sky130_fd_sc_hd__nor2_1 _06290_ (.A(_00443_),
    .B(_00444_),
    .Y(_00445_));
 sky130_fd_sc_hd__xor2_1 _06291_ (.A(_00443_),
    .B(_00444_),
    .X(_00446_));
 sky130_fd_sc_hd__xor2_1 _06292_ (.A(_00325_),
    .B(_00446_),
    .X(_00447_));
 sky130_fd_sc_hd__and3_1 _06293_ (.A(net1),
    .B(net48),
    .C(_00447_),
    .X(_00448_));
 sky130_fd_sc_hd__a21oi_1 _06294_ (.A1(net1),
    .A2(net48),
    .B1(_00447_),
    .Y(_00449_));
 sky130_fd_sc_hd__nor2_1 _06295_ (.A(_00448_),
    .B(_00449_),
    .Y(\genblk2[22].rca.ripple_adders[23].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _06296_ (.A1(_00325_),
    .A2(_00446_),
    .B1(_00445_),
    .X(_00451_));
 sky130_fd_sc_hd__a21o_1 _06297_ (.A1(_00327_),
    .A2(_00442_),
    .B1(_00441_),
    .X(_00452_));
 sky130_fd_sc_hd__a21o_1 _06298_ (.A1(_00328_),
    .A2(_00437_),
    .B1(_00436_),
    .X(_00453_));
 sky130_fd_sc_hd__a21o_1 _06299_ (.A1(_00330_),
    .A2(_00433_),
    .B1(_00432_),
    .X(_00454_));
 sky130_fd_sc_hd__a21o_1 _06300_ (.A1(_00331_),
    .A2(_00429_),
    .B1(_00427_),
    .X(_00455_));
 sky130_fd_sc_hd__a21o_1 _06301_ (.A1(_00332_),
    .A2(_00424_),
    .B1(_00423_),
    .X(_00456_));
 sky130_fd_sc_hd__a21o_1 _06302_ (.A1(_00333_),
    .A2(_00420_),
    .B1(_00419_),
    .X(_00457_));
 sky130_fd_sc_hd__a21o_1 _06303_ (.A1(_00334_),
    .A2(_00415_),
    .B1(_00414_),
    .X(_00458_));
 sky130_fd_sc_hd__a21o_1 _06304_ (.A1(_00335_),
    .A2(_00411_),
    .B1(_00410_),
    .X(_00459_));
 sky130_fd_sc_hd__a21o_1 _06305_ (.A1(_00336_),
    .A2(_00407_),
    .B1(_00405_),
    .X(_00461_));
 sky130_fd_sc_hd__a21o_1 _06306_ (.A1(_00337_),
    .A2(_00402_),
    .B1(_00401_),
    .X(_00462_));
 sky130_fd_sc_hd__a21o_1 _06307_ (.A1(_00338_),
    .A2(_00398_),
    .B1(_00397_),
    .X(_00463_));
 sky130_fd_sc_hd__a21o_1 _06308_ (.A1(_00339_),
    .A2(_00393_),
    .B1(_00392_),
    .X(_00464_));
 sky130_fd_sc_hd__a21o_1 _06309_ (.A1(_00341_),
    .A2(_00389_),
    .B1(_00388_),
    .X(_00465_));
 sky130_fd_sc_hd__a21o_1 _06310_ (.A1(_00342_),
    .A2(_00385_),
    .B1(_00383_),
    .X(_00466_));
 sky130_fd_sc_hd__a21o_1 _06311_ (.A1(_00343_),
    .A2(_00380_),
    .B1(_00379_),
    .X(_00467_));
 sky130_fd_sc_hd__a21o_1 _06312_ (.A1(_00344_),
    .A2(_00376_),
    .B1(_00375_),
    .X(_00468_));
 sky130_fd_sc_hd__a21o_1 _06313_ (.A1(_00345_),
    .A2(_00371_),
    .B1(_00370_),
    .X(_00469_));
 sky130_fd_sc_hd__a21o_1 _06314_ (.A1(_00346_),
    .A2(_00367_),
    .B1(_00366_),
    .X(_00470_));
 sky130_fd_sc_hd__a21o_1 _06315_ (.A1(_00347_),
    .A2(_00363_),
    .B1(_00361_),
    .X(_00472_));
 sky130_fd_sc_hd__a21o_1 _06316_ (.A1(_00348_),
    .A2(_00357_),
    .B1(_00356_),
    .X(_00473_));
 sky130_fd_sc_hd__a22o_1 _06317_ (.A1(net44),
    .A2(net16),
    .B1(net17),
    .B2(net33),
    .X(_00474_));
 sky130_fd_sc_hd__and3_1 _06318_ (.A(net44),
    .B(net16),
    .C(net17),
    .X(_00475_));
 sky130_fd_sc_hd__a21bo_1 _06319_ (.A1(net33),
    .A2(_00475_),
    .B1_N(_00474_),
    .X(_00476_));
 sky130_fd_sc_hd__a22o_1 _06320_ (.A1(net33),
    .A2(_00350_),
    .B1(_00353_),
    .B2(_00349_),
    .X(_00477_));
 sky130_fd_sc_hd__xnor2_1 _06321_ (.A(_00476_),
    .B(_00477_),
    .Y(_00478_));
 sky130_fd_sc_hd__nand2_1 _06322_ (.A(net55),
    .B(net15),
    .Y(_00479_));
 sky130_fd_sc_hd__and3_1 _06323_ (.A(net55),
    .B(net15),
    .C(_00478_),
    .X(_00480_));
 sky130_fd_sc_hd__nand2b_1 _06324_ (.A_N(_00478_),
    .B(_00479_),
    .Y(_00481_));
 sky130_fd_sc_hd__xor2_1 _06325_ (.A(_00478_),
    .B(_00479_),
    .X(_00483_));
 sky130_fd_sc_hd__xnor2_1 _06326_ (.A(_00473_),
    .B(_00483_),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_1 _06327_ (.A(net58),
    .B(net14),
    .Y(_00485_));
 sky130_fd_sc_hd__and3_1 _06328_ (.A(net58),
    .B(net14),
    .C(_00484_),
    .X(_00486_));
 sky130_fd_sc_hd__xnor2_1 _06329_ (.A(_00484_),
    .B(_00485_),
    .Y(_00487_));
 sky130_fd_sc_hd__xor2_1 _06330_ (.A(_00472_),
    .B(_00487_),
    .X(_00488_));
 sky130_fd_sc_hd__nand2_1 _06331_ (.A(net59),
    .B(net13),
    .Y(_00489_));
 sky130_fd_sc_hd__and3_1 _06332_ (.A(net59),
    .B(net13),
    .C(_00488_),
    .X(_00490_));
 sky130_fd_sc_hd__xnor2_1 _06333_ (.A(_00488_),
    .B(_00489_),
    .Y(_00491_));
 sky130_fd_sc_hd__xor2_1 _06334_ (.A(_00470_),
    .B(_00491_),
    .X(_00492_));
 sky130_fd_sc_hd__nand2_1 _06335_ (.A(net60),
    .B(net11),
    .Y(_00494_));
 sky130_fd_sc_hd__and3_1 _06336_ (.A(net60),
    .B(net11),
    .C(_00492_),
    .X(_00495_));
 sky130_fd_sc_hd__xnor2_1 _06337_ (.A(_00492_),
    .B(_00494_),
    .Y(_00496_));
 sky130_fd_sc_hd__xor2_1 _06338_ (.A(_00469_),
    .B(_00496_),
    .X(_00497_));
 sky130_fd_sc_hd__nand2_1 _06339_ (.A(net61),
    .B(net10),
    .Y(_00498_));
 sky130_fd_sc_hd__and3_1 _06340_ (.A(net61),
    .B(net10),
    .C(_00497_),
    .X(_00499_));
 sky130_fd_sc_hd__xnor2_1 _06341_ (.A(_00497_),
    .B(_00498_),
    .Y(_00500_));
 sky130_fd_sc_hd__xor2_1 _06342_ (.A(_00468_),
    .B(_00500_),
    .X(_00501_));
 sky130_fd_sc_hd__nand2_1 _06343_ (.A(net62),
    .B(net9),
    .Y(_00502_));
 sky130_fd_sc_hd__and3_1 _06344_ (.A(net62),
    .B(net9),
    .C(_00501_),
    .X(_00503_));
 sky130_fd_sc_hd__xnor2_1 _06345_ (.A(_00501_),
    .B(_00502_),
    .Y(_00505_));
 sky130_fd_sc_hd__xnor2_1 _06346_ (.A(_00467_),
    .B(_00505_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_1 _06347_ (.A(net63),
    .B(net8),
    .Y(_00507_));
 sky130_fd_sc_hd__nor2_1 _06348_ (.A(_00506_),
    .B(_00507_),
    .Y(_00508_));
 sky130_fd_sc_hd__xor2_1 _06349_ (.A(_00506_),
    .B(_00507_),
    .X(_00509_));
 sky130_fd_sc_hd__xnor2_1 _06350_ (.A(_00466_),
    .B(_00509_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _06351_ (.A(net64),
    .B(net7),
    .Y(_00511_));
 sky130_fd_sc_hd__nor2_1 _06352_ (.A(_00510_),
    .B(_00511_),
    .Y(_00512_));
 sky130_fd_sc_hd__xor2_1 _06353_ (.A(_00510_),
    .B(_00511_),
    .X(_00513_));
 sky130_fd_sc_hd__xnor2_1 _06354_ (.A(_00465_),
    .B(_00513_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand2_1 _06355_ (.A(net34),
    .B(net6),
    .Y(_00516_));
 sky130_fd_sc_hd__nor2_1 _06356_ (.A(_00514_),
    .B(_00516_),
    .Y(_00517_));
 sky130_fd_sc_hd__xor2_1 _06357_ (.A(_00514_),
    .B(_00516_),
    .X(_00518_));
 sky130_fd_sc_hd__xnor2_1 _06358_ (.A(_00464_),
    .B(_00518_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_1 _06359_ (.A(net35),
    .B(net5),
    .Y(_00520_));
 sky130_fd_sc_hd__nor2_1 _06360_ (.A(_00519_),
    .B(_00520_),
    .Y(_00521_));
 sky130_fd_sc_hd__xor2_1 _06361_ (.A(_00519_),
    .B(_00520_),
    .X(_00522_));
 sky130_fd_sc_hd__xnor2_1 _06362_ (.A(_00463_),
    .B(_00522_),
    .Y(_00523_));
 sky130_fd_sc_hd__nand2_1 _06363_ (.A(net36),
    .B(net4),
    .Y(_00524_));
 sky130_fd_sc_hd__nor2_1 _06364_ (.A(_00523_),
    .B(_00524_),
    .Y(_00525_));
 sky130_fd_sc_hd__xor2_1 _06365_ (.A(_00523_),
    .B(_00524_),
    .X(_00527_));
 sky130_fd_sc_hd__xnor2_1 _06366_ (.A(_00462_),
    .B(_00527_),
    .Y(_00528_));
 sky130_fd_sc_hd__nand2_1 _06367_ (.A(net3),
    .B(net37),
    .Y(_00529_));
 sky130_fd_sc_hd__nor2_1 _06368_ (.A(_00528_),
    .B(_00529_),
    .Y(_00530_));
 sky130_fd_sc_hd__xor2_1 _06369_ (.A(_00528_),
    .B(_00529_),
    .X(_00531_));
 sky130_fd_sc_hd__xnor2_1 _06370_ (.A(_00461_),
    .B(_00531_),
    .Y(_00532_));
 sky130_fd_sc_hd__nand2_1 _06371_ (.A(net2),
    .B(net38),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2_1 _06372_ (.A(_00532_),
    .B(_00533_),
    .Y(_00534_));
 sky130_fd_sc_hd__xor2_1 _06373_ (.A(_00532_),
    .B(_00533_),
    .X(_00535_));
 sky130_fd_sc_hd__xnor2_1 _06374_ (.A(_00459_),
    .B(_00535_),
    .Y(_00536_));
 sky130_fd_sc_hd__nand2_1 _06375_ (.A(net32),
    .B(net39),
    .Y(_00538_));
 sky130_fd_sc_hd__nor2_1 _06376_ (.A(_00536_),
    .B(_00538_),
    .Y(_00539_));
 sky130_fd_sc_hd__xor2_1 _06377_ (.A(_00536_),
    .B(_00538_),
    .X(_00540_));
 sky130_fd_sc_hd__xnor2_1 _06378_ (.A(_00458_),
    .B(_00540_),
    .Y(_00541_));
 sky130_fd_sc_hd__nand2_1 _06379_ (.A(net31),
    .B(net40),
    .Y(_00542_));
 sky130_fd_sc_hd__nor2_1 _06380_ (.A(_00541_),
    .B(_00542_),
    .Y(_00543_));
 sky130_fd_sc_hd__xor2_1 _06381_ (.A(_00541_),
    .B(_00542_),
    .X(_00544_));
 sky130_fd_sc_hd__xnor2_1 _06382_ (.A(_00457_),
    .B(_00544_),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2_1 _06383_ (.A(net30),
    .B(net41),
    .Y(_00546_));
 sky130_fd_sc_hd__nor2_1 _06384_ (.A(_00545_),
    .B(_00546_),
    .Y(_00547_));
 sky130_fd_sc_hd__xor2_1 _06385_ (.A(_00545_),
    .B(_00546_),
    .X(_00549_));
 sky130_fd_sc_hd__xnor2_1 _06386_ (.A(_00456_),
    .B(_00549_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2_1 _06387_ (.A(net29),
    .B(net42),
    .Y(_00551_));
 sky130_fd_sc_hd__nor2_1 _06388_ (.A(_00550_),
    .B(_00551_),
    .Y(_00552_));
 sky130_fd_sc_hd__xor2_1 _06389_ (.A(_00550_),
    .B(_00551_),
    .X(_00553_));
 sky130_fd_sc_hd__xnor2_1 _06390_ (.A(_00455_),
    .B(_00553_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2_1 _06391_ (.A(net28),
    .B(net43),
    .Y(_00555_));
 sky130_fd_sc_hd__nor2_1 _06392_ (.A(_00554_),
    .B(_00555_),
    .Y(_00556_));
 sky130_fd_sc_hd__xor2_1 _06393_ (.A(_00554_),
    .B(_00555_),
    .X(_00557_));
 sky130_fd_sc_hd__xnor2_1 _06394_ (.A(_00454_),
    .B(_00557_),
    .Y(_00558_));
 sky130_fd_sc_hd__nand2_1 _06395_ (.A(net27),
    .B(net45),
    .Y(_00560_));
 sky130_fd_sc_hd__nor2_1 _06396_ (.A(_00558_),
    .B(_00560_),
    .Y(_00561_));
 sky130_fd_sc_hd__xor2_1 _06397_ (.A(_00558_),
    .B(_00560_),
    .X(_00562_));
 sky130_fd_sc_hd__xnor2_1 _06398_ (.A(_00453_),
    .B(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand2_1 _06399_ (.A(net26),
    .B(net46),
    .Y(_00564_));
 sky130_fd_sc_hd__nor2_1 _06400_ (.A(_00563_),
    .B(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__xor2_1 _06401_ (.A(_00563_),
    .B(_00564_),
    .X(_00566_));
 sky130_fd_sc_hd__xnor2_1 _06402_ (.A(_00452_),
    .B(_00566_),
    .Y(_00567_));
 sky130_fd_sc_hd__nand2_1 _06403_ (.A(net23),
    .B(net47),
    .Y(_00568_));
 sky130_fd_sc_hd__nor2_1 _06404_ (.A(_00567_),
    .B(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__xor2_1 _06405_ (.A(_00567_),
    .B(_00568_),
    .X(_00571_));
 sky130_fd_sc_hd__xnor2_1 _06406_ (.A(_00451_),
    .B(_00571_),
    .Y(_00572_));
 sky130_fd_sc_hd__nand2_1 _06407_ (.A(net12),
    .B(net48),
    .Y(_00573_));
 sky130_fd_sc_hd__nor2_1 _06408_ (.A(_00572_),
    .B(_00573_),
    .Y(_00574_));
 sky130_fd_sc_hd__xor2_1 _06409_ (.A(_00572_),
    .B(_00573_),
    .X(_00575_));
 sky130_fd_sc_hd__xor2_1 _06410_ (.A(_00448_),
    .B(_00575_),
    .X(_00576_));
 sky130_fd_sc_hd__and3_1 _06411_ (.A(net1),
    .B(net49),
    .C(_00576_),
    .X(_00577_));
 sky130_fd_sc_hd__a21oi_1 _06412_ (.A1(net1),
    .A2(net49),
    .B1(_00576_),
    .Y(_00578_));
 sky130_fd_sc_hd__nor2_1 _06413_ (.A(_00577_),
    .B(_00578_),
    .Y(\genblk2[23].rca.ripple_adders[24].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _06414_ (.A1(_00448_),
    .A2(_00575_),
    .B1(_00574_),
    .X(_00579_));
 sky130_fd_sc_hd__a21o_1 _06415_ (.A1(_00451_),
    .A2(_00571_),
    .B1(_00569_),
    .X(_00581_));
 sky130_fd_sc_hd__a21o_1 _06416_ (.A1(_00452_),
    .A2(_00566_),
    .B1(_00565_),
    .X(_00582_));
 sky130_fd_sc_hd__a21o_1 _06417_ (.A1(_00453_),
    .A2(_00562_),
    .B1(_00561_),
    .X(_00583_));
 sky130_fd_sc_hd__a21o_1 _06418_ (.A1(_00454_),
    .A2(_00557_),
    .B1(_00556_),
    .X(_00584_));
 sky130_fd_sc_hd__a21o_1 _06419_ (.A1(_00455_),
    .A2(_00553_),
    .B1(_00552_),
    .X(_00585_));
 sky130_fd_sc_hd__a21o_1 _06420_ (.A1(_00456_),
    .A2(_00549_),
    .B1(_00547_),
    .X(_00586_));
 sky130_fd_sc_hd__a21o_1 _06421_ (.A1(_00457_),
    .A2(_00544_),
    .B1(_00543_),
    .X(_00587_));
 sky130_fd_sc_hd__a21o_1 _06422_ (.A1(_00458_),
    .A2(_00540_),
    .B1(_00539_),
    .X(_00588_));
 sky130_fd_sc_hd__a21o_1 _06423_ (.A1(_00459_),
    .A2(_00535_),
    .B1(_00534_),
    .X(_00589_));
 sky130_fd_sc_hd__a21o_1 _06424_ (.A1(_00461_),
    .A2(_00531_),
    .B1(_00530_),
    .X(_00590_));
 sky130_fd_sc_hd__a21o_1 _06425_ (.A1(_00462_),
    .A2(_00527_),
    .B1(_00525_),
    .X(_00592_));
 sky130_fd_sc_hd__a21o_1 _06426_ (.A1(_00463_),
    .A2(_00522_),
    .B1(_00521_),
    .X(_00593_));
 sky130_fd_sc_hd__a21o_1 _06427_ (.A1(_00464_),
    .A2(_00518_),
    .B1(_00517_),
    .X(_00594_));
 sky130_fd_sc_hd__a21o_1 _06428_ (.A1(_00465_),
    .A2(_00513_),
    .B1(_00512_),
    .X(_00595_));
 sky130_fd_sc_hd__a21o_1 _06429_ (.A1(_00466_),
    .A2(_00509_),
    .B1(_00508_),
    .X(_00596_));
 sky130_fd_sc_hd__a21o_1 _06430_ (.A1(_00467_),
    .A2(_00505_),
    .B1(_00503_),
    .X(_00597_));
 sky130_fd_sc_hd__a21o_1 _06431_ (.A1(_00468_),
    .A2(_00500_),
    .B1(_00499_),
    .X(_00598_));
 sky130_fd_sc_hd__a21o_1 _06432_ (.A1(_00469_),
    .A2(_00496_),
    .B1(_00495_),
    .X(_00599_));
 sky130_fd_sc_hd__a21o_1 _06433_ (.A1(_00470_),
    .A2(_00491_),
    .B1(_00490_),
    .X(_00600_));
 sky130_fd_sc_hd__a21o_1 _06434_ (.A1(_00472_),
    .A2(_00487_),
    .B1(_00486_),
    .X(_00601_));
 sky130_fd_sc_hd__a21o_1 _06435_ (.A1(_00473_),
    .A2(_00481_),
    .B1(_00480_),
    .X(_00603_));
 sky130_fd_sc_hd__a22o_1 _06436_ (.A1(net44),
    .A2(net17),
    .B1(net18),
    .B2(net33),
    .X(_00604_));
 sky130_fd_sc_hd__and3_1 _06437_ (.A(net44),
    .B(net17),
    .C(net18),
    .X(_00605_));
 sky130_fd_sc_hd__a21bo_1 _06438_ (.A1(net33),
    .A2(_00605_),
    .B1_N(_00604_),
    .X(_00606_));
 sky130_fd_sc_hd__a22o_1 _06439_ (.A1(net33),
    .A2(_00475_),
    .B1(_00477_),
    .B2(_00474_),
    .X(_00607_));
 sky130_fd_sc_hd__xnor2_1 _06440_ (.A(_00606_),
    .B(_00607_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _06441_ (.A(net55),
    .B(net16),
    .Y(_00609_));
 sky130_fd_sc_hd__and3_1 _06442_ (.A(net55),
    .B(net16),
    .C(_00608_),
    .X(_00610_));
 sky130_fd_sc_hd__nand2b_1 _06443_ (.A_N(_00608_),
    .B(_00609_),
    .Y(_00611_));
 sky130_fd_sc_hd__xor2_1 _06444_ (.A(_00608_),
    .B(_00609_),
    .X(_00612_));
 sky130_fd_sc_hd__xnor2_1 _06445_ (.A(_00603_),
    .B(_00612_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_1 _06446_ (.A(net58),
    .B(net15),
    .Y(_00615_));
 sky130_fd_sc_hd__and3_1 _06447_ (.A(net58),
    .B(net15),
    .C(_00614_),
    .X(_00616_));
 sky130_fd_sc_hd__xnor2_1 _06448_ (.A(_00614_),
    .B(_00615_),
    .Y(_00617_));
 sky130_fd_sc_hd__xor2_1 _06449_ (.A(_00601_),
    .B(_00617_),
    .X(_00618_));
 sky130_fd_sc_hd__nand2_1 _06450_ (.A(net59),
    .B(net14),
    .Y(_00619_));
 sky130_fd_sc_hd__and3_1 _06451_ (.A(net59),
    .B(net14),
    .C(_00618_),
    .X(_00620_));
 sky130_fd_sc_hd__xnor2_1 _06452_ (.A(_00618_),
    .B(_00619_),
    .Y(_00621_));
 sky130_fd_sc_hd__xor2_1 _06453_ (.A(_00600_),
    .B(_00621_),
    .X(_00622_));
 sky130_fd_sc_hd__nand2_1 _06454_ (.A(net60),
    .B(net13),
    .Y(_00623_));
 sky130_fd_sc_hd__and3_1 _06455_ (.A(net60),
    .B(net13),
    .C(_00622_),
    .X(_00625_));
 sky130_fd_sc_hd__xnor2_1 _06456_ (.A(_00622_),
    .B(_00623_),
    .Y(_00626_));
 sky130_fd_sc_hd__xor2_1 _06457_ (.A(_00599_),
    .B(_00626_),
    .X(_00627_));
 sky130_fd_sc_hd__nand2_1 _06458_ (.A(net61),
    .B(net11),
    .Y(_00628_));
 sky130_fd_sc_hd__and3_1 _06459_ (.A(net61),
    .B(net11),
    .C(_00627_),
    .X(_00629_));
 sky130_fd_sc_hd__xnor2_1 _06460_ (.A(_00627_),
    .B(_00628_),
    .Y(_00630_));
 sky130_fd_sc_hd__xor2_1 _06461_ (.A(_00598_),
    .B(_00630_),
    .X(_00631_));
 sky130_fd_sc_hd__nand2_1 _06462_ (.A(net62),
    .B(net10),
    .Y(_00632_));
 sky130_fd_sc_hd__and3_1 _06463_ (.A(net62),
    .B(net10),
    .C(_00631_),
    .X(_00633_));
 sky130_fd_sc_hd__xnor2_1 _06464_ (.A(_00631_),
    .B(_00632_),
    .Y(_00634_));
 sky130_fd_sc_hd__xnor2_1 _06465_ (.A(_00597_),
    .B(_00634_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _06466_ (.A(net63),
    .B(net9),
    .Y(_00637_));
 sky130_fd_sc_hd__nor2_1 _06467_ (.A(_00636_),
    .B(_00637_),
    .Y(_00638_));
 sky130_fd_sc_hd__xor2_1 _06468_ (.A(_00636_),
    .B(_00637_),
    .X(_00639_));
 sky130_fd_sc_hd__xnor2_1 _06469_ (.A(_00596_),
    .B(_00639_),
    .Y(_00640_));
 sky130_fd_sc_hd__nand2_1 _06470_ (.A(net64),
    .B(net8),
    .Y(_00641_));
 sky130_fd_sc_hd__nor2_1 _06471_ (.A(_00640_),
    .B(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hd__xor2_1 _06472_ (.A(_00640_),
    .B(_00641_),
    .X(_00643_));
 sky130_fd_sc_hd__xnor2_1 _06473_ (.A(_00595_),
    .B(_00643_),
    .Y(_00644_));
 sky130_fd_sc_hd__nand2_1 _06474_ (.A(net34),
    .B(net7),
    .Y(_00645_));
 sky130_fd_sc_hd__nor2_1 _06475_ (.A(_00644_),
    .B(_00645_),
    .Y(_00647_));
 sky130_fd_sc_hd__xor2_1 _06476_ (.A(_00644_),
    .B(_00645_),
    .X(_00648_));
 sky130_fd_sc_hd__xnor2_1 _06477_ (.A(_00594_),
    .B(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__nand2_1 _06478_ (.A(net35),
    .B(net6),
    .Y(_00650_));
 sky130_fd_sc_hd__nor2_1 _06479_ (.A(_00649_),
    .B(_00650_),
    .Y(_00651_));
 sky130_fd_sc_hd__xor2_1 _06480_ (.A(_00649_),
    .B(_00650_),
    .X(_00652_));
 sky130_fd_sc_hd__xnor2_1 _06481_ (.A(_00593_),
    .B(_00652_),
    .Y(_00653_));
 sky130_fd_sc_hd__nand2_1 _06482_ (.A(net36),
    .B(net5),
    .Y(_00654_));
 sky130_fd_sc_hd__nor2_1 _06483_ (.A(_00653_),
    .B(_00654_),
    .Y(_00655_));
 sky130_fd_sc_hd__xor2_1 _06484_ (.A(_00653_),
    .B(_00654_),
    .X(_00656_));
 sky130_fd_sc_hd__xnor2_1 _06485_ (.A(_00592_),
    .B(_00656_),
    .Y(_00658_));
 sky130_fd_sc_hd__nand2_1 _06486_ (.A(net4),
    .B(net37),
    .Y(_00659_));
 sky130_fd_sc_hd__nor2_1 _06487_ (.A(_00658_),
    .B(_00659_),
    .Y(_00660_));
 sky130_fd_sc_hd__xor2_1 _06488_ (.A(_00658_),
    .B(_00659_),
    .X(_00661_));
 sky130_fd_sc_hd__xnor2_1 _06489_ (.A(_00590_),
    .B(_00661_),
    .Y(_00662_));
 sky130_fd_sc_hd__nand2_1 _06490_ (.A(net3),
    .B(net38),
    .Y(_00663_));
 sky130_fd_sc_hd__nor2_1 _06491_ (.A(_00662_),
    .B(_00663_),
    .Y(_00664_));
 sky130_fd_sc_hd__xor2_1 _06492_ (.A(_00662_),
    .B(_00663_),
    .X(_00665_));
 sky130_fd_sc_hd__xnor2_1 _06493_ (.A(_00589_),
    .B(_00665_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_1 _06494_ (.A(net2),
    .B(net39),
    .Y(_00667_));
 sky130_fd_sc_hd__nor2_1 _06495_ (.A(_00666_),
    .B(_00667_),
    .Y(_00669_));
 sky130_fd_sc_hd__xor2_1 _06496_ (.A(_00666_),
    .B(_00667_),
    .X(_00670_));
 sky130_fd_sc_hd__xnor2_1 _06497_ (.A(_00588_),
    .B(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__nand2_1 _06498_ (.A(net32),
    .B(net40),
    .Y(_00672_));
 sky130_fd_sc_hd__nor2_1 _06499_ (.A(_00671_),
    .B(_00672_),
    .Y(_00673_));
 sky130_fd_sc_hd__xor2_1 _06500_ (.A(_00671_),
    .B(_00672_),
    .X(_00674_));
 sky130_fd_sc_hd__xnor2_1 _06501_ (.A(_00587_),
    .B(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__nand2_1 _06502_ (.A(net31),
    .B(net41),
    .Y(_00676_));
 sky130_fd_sc_hd__nor2_1 _06503_ (.A(_00675_),
    .B(_00676_),
    .Y(_00677_));
 sky130_fd_sc_hd__xor2_1 _06504_ (.A(_00675_),
    .B(_00676_),
    .X(_00678_));
 sky130_fd_sc_hd__xnor2_1 _06505_ (.A(_00586_),
    .B(_00678_),
    .Y(_00680_));
 sky130_fd_sc_hd__nand2_1 _06506_ (.A(net30),
    .B(net42),
    .Y(_00681_));
 sky130_fd_sc_hd__nor2_1 _06507_ (.A(_00680_),
    .B(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__xor2_1 _06508_ (.A(_00680_),
    .B(_00681_),
    .X(_00683_));
 sky130_fd_sc_hd__xnor2_1 _06509_ (.A(_00585_),
    .B(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__nand2_1 _06510_ (.A(net29),
    .B(net43),
    .Y(_00685_));
 sky130_fd_sc_hd__nor2_1 _06511_ (.A(_00684_),
    .B(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__xor2_1 _06512_ (.A(_00684_),
    .B(_00685_),
    .X(_00687_));
 sky130_fd_sc_hd__xnor2_1 _06513_ (.A(_00584_),
    .B(_00687_),
    .Y(_00688_));
 sky130_fd_sc_hd__nand2_1 _06514_ (.A(net28),
    .B(net45),
    .Y(_00689_));
 sky130_fd_sc_hd__nor2_1 _06515_ (.A(_00688_),
    .B(_00689_),
    .Y(_00691_));
 sky130_fd_sc_hd__xor2_1 _06516_ (.A(_00688_),
    .B(_00689_),
    .X(_00692_));
 sky130_fd_sc_hd__xnor2_1 _06517_ (.A(_00583_),
    .B(_00692_),
    .Y(_00693_));
 sky130_fd_sc_hd__nand2_1 _06518_ (.A(net27),
    .B(net46),
    .Y(_00694_));
 sky130_fd_sc_hd__nor2_1 _06519_ (.A(_00693_),
    .B(_00694_),
    .Y(_00695_));
 sky130_fd_sc_hd__xor2_1 _06520_ (.A(_00693_),
    .B(_00694_),
    .X(_00696_));
 sky130_fd_sc_hd__xnor2_1 _06521_ (.A(_00582_),
    .B(_00696_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand2_1 _06522_ (.A(net26),
    .B(net47),
    .Y(_00698_));
 sky130_fd_sc_hd__nor2_1 _06523_ (.A(_00697_),
    .B(_00698_),
    .Y(_00699_));
 sky130_fd_sc_hd__xor2_1 _06524_ (.A(_00697_),
    .B(_00698_),
    .X(_00700_));
 sky130_fd_sc_hd__xnor2_1 _06525_ (.A(_00581_),
    .B(_00700_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand2_1 _06526_ (.A(net23),
    .B(net48),
    .Y(_00703_));
 sky130_fd_sc_hd__nor2_1 _06527_ (.A(_00702_),
    .B(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__xor2_1 _06528_ (.A(_00702_),
    .B(_00703_),
    .X(_00705_));
 sky130_fd_sc_hd__xnor2_1 _06529_ (.A(_00579_),
    .B(_00705_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand2_1 _06530_ (.A(net12),
    .B(net49),
    .Y(_00707_));
 sky130_fd_sc_hd__nor2_1 _06531_ (.A(_00706_),
    .B(_00707_),
    .Y(_00708_));
 sky130_fd_sc_hd__xor2_1 _06532_ (.A(_00706_),
    .B(_00707_),
    .X(_00709_));
 sky130_fd_sc_hd__xor2_1 _06533_ (.A(_00577_),
    .B(_00709_),
    .X(_00710_));
 sky130_fd_sc_hd__and3_1 _06534_ (.A(net1),
    .B(net50),
    .C(_00710_),
    .X(_00711_));
 sky130_fd_sc_hd__a21oi_1 _06535_ (.A1(net1),
    .A2(net50),
    .B1(_00710_),
    .Y(_00713_));
 sky130_fd_sc_hd__nor2_1 _06536_ (.A(_00711_),
    .B(_00713_),
    .Y(\genblk2[24].rca.ripple_adders[25].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _06537_ (.A1(_00577_),
    .A2(_00709_),
    .B1(_00708_),
    .X(_00714_));
 sky130_fd_sc_hd__a21o_1 _06538_ (.A1(_00579_),
    .A2(_00705_),
    .B1(_00704_),
    .X(_00715_));
 sky130_fd_sc_hd__a21o_1 _06539_ (.A1(_00581_),
    .A2(_00700_),
    .B1(_00699_),
    .X(_00716_));
 sky130_fd_sc_hd__a21o_1 _06540_ (.A1(_00582_),
    .A2(_00696_),
    .B1(_00695_),
    .X(_00717_));
 sky130_fd_sc_hd__a21o_1 _06541_ (.A1(_00583_),
    .A2(_00692_),
    .B1(_00691_),
    .X(_00718_));
 sky130_fd_sc_hd__a21o_1 _06542_ (.A1(_00584_),
    .A2(_00687_),
    .B1(_00686_),
    .X(_00719_));
 sky130_fd_sc_hd__a21o_1 _06543_ (.A1(_00585_),
    .A2(_00683_),
    .B1(_00682_),
    .X(_00720_));
 sky130_fd_sc_hd__a21o_1 _06544_ (.A1(_00586_),
    .A2(_00678_),
    .B1(_00677_),
    .X(_00721_));
 sky130_fd_sc_hd__a21o_1 _06545_ (.A1(_00587_),
    .A2(_00674_),
    .B1(_00673_),
    .X(_00723_));
 sky130_fd_sc_hd__a21o_1 _06546_ (.A1(_00588_),
    .A2(_00670_),
    .B1(_00669_),
    .X(_00724_));
 sky130_fd_sc_hd__a21o_1 _06547_ (.A1(_00589_),
    .A2(_00665_),
    .B1(_00664_),
    .X(_00725_));
 sky130_fd_sc_hd__a21o_1 _06548_ (.A1(_00590_),
    .A2(_00661_),
    .B1(_00660_),
    .X(_00726_));
 sky130_fd_sc_hd__a21o_1 _06549_ (.A1(_00592_),
    .A2(_00656_),
    .B1(_00655_),
    .X(_00727_));
 sky130_fd_sc_hd__a21o_1 _06550_ (.A1(_00593_),
    .A2(_00652_),
    .B1(_00651_),
    .X(_00728_));
 sky130_fd_sc_hd__a21o_1 _06551_ (.A1(_00594_),
    .A2(_00648_),
    .B1(_00647_),
    .X(_00729_));
 sky130_fd_sc_hd__a21o_1 _06552_ (.A1(_00595_),
    .A2(_00643_),
    .B1(_00642_),
    .X(_00730_));
 sky130_fd_sc_hd__a21o_1 _06553_ (.A1(_00596_),
    .A2(_00639_),
    .B1(_00638_),
    .X(_00731_));
 sky130_fd_sc_hd__a21o_1 _06554_ (.A1(_00597_),
    .A2(_00634_),
    .B1(_00633_),
    .X(_00732_));
 sky130_fd_sc_hd__a21o_1 _06555_ (.A1(_00598_),
    .A2(_00630_),
    .B1(_00629_),
    .X(_00734_));
 sky130_fd_sc_hd__a21o_1 _06556_ (.A1(_00599_),
    .A2(_00626_),
    .B1(_00625_),
    .X(_00735_));
 sky130_fd_sc_hd__a21o_1 _06557_ (.A1(_00600_),
    .A2(_00621_),
    .B1(_00620_),
    .X(_00736_));
 sky130_fd_sc_hd__a21o_1 _06558_ (.A1(_00601_),
    .A2(_00617_),
    .B1(_00616_),
    .X(_00737_));
 sky130_fd_sc_hd__a21o_1 _06559_ (.A1(_00603_),
    .A2(_00611_),
    .B1(_00610_),
    .X(_00738_));
 sky130_fd_sc_hd__a22o_1 _06560_ (.A1(net44),
    .A2(net18),
    .B1(net19),
    .B2(net33),
    .X(_00739_));
 sky130_fd_sc_hd__and3_1 _06561_ (.A(net44),
    .B(net18),
    .C(net19),
    .X(_00740_));
 sky130_fd_sc_hd__a21bo_1 _06562_ (.A1(net33),
    .A2(_00740_),
    .B1_N(_00739_),
    .X(_00741_));
 sky130_fd_sc_hd__a22o_1 _06563_ (.A1(net33),
    .A2(_00605_),
    .B1(_00607_),
    .B2(_00604_),
    .X(_00742_));
 sky130_fd_sc_hd__xnor2_1 _06564_ (.A(_00741_),
    .B(_00742_),
    .Y(_00743_));
 sky130_fd_sc_hd__nand2_1 _06565_ (.A(net55),
    .B(net17),
    .Y(_00745_));
 sky130_fd_sc_hd__and3_1 _06566_ (.A(net55),
    .B(net17),
    .C(_00743_),
    .X(_00746_));
 sky130_fd_sc_hd__nand2b_1 _06567_ (.A_N(_00743_),
    .B(_00745_),
    .Y(_00747_));
 sky130_fd_sc_hd__xor2_1 _06568_ (.A(_00743_),
    .B(_00745_),
    .X(_00748_));
 sky130_fd_sc_hd__xnor2_1 _06569_ (.A(_00738_),
    .B(_00748_),
    .Y(_00749_));
 sky130_fd_sc_hd__nand2_1 _06570_ (.A(net58),
    .B(net16),
    .Y(_00750_));
 sky130_fd_sc_hd__and3_1 _06571_ (.A(net58),
    .B(net16),
    .C(_00749_),
    .X(_00751_));
 sky130_fd_sc_hd__xnor2_1 _06572_ (.A(_00749_),
    .B(_00750_),
    .Y(_00752_));
 sky130_fd_sc_hd__xor2_1 _06573_ (.A(_00737_),
    .B(_00752_),
    .X(_00753_));
 sky130_fd_sc_hd__nand2_1 _06574_ (.A(net59),
    .B(net15),
    .Y(_00754_));
 sky130_fd_sc_hd__and3_1 _06575_ (.A(net59),
    .B(net15),
    .C(_00753_),
    .X(_00756_));
 sky130_fd_sc_hd__xnor2_1 _06576_ (.A(_00753_),
    .B(_00754_),
    .Y(_00757_));
 sky130_fd_sc_hd__xor2_1 _06577_ (.A(_00736_),
    .B(_00757_),
    .X(_00758_));
 sky130_fd_sc_hd__nand2_1 _06578_ (.A(net60),
    .B(net14),
    .Y(_00759_));
 sky130_fd_sc_hd__and3_1 _06579_ (.A(net60),
    .B(net14),
    .C(_00758_),
    .X(_00760_));
 sky130_fd_sc_hd__xnor2_1 _06580_ (.A(_00758_),
    .B(_00759_),
    .Y(_00761_));
 sky130_fd_sc_hd__xor2_1 _06581_ (.A(_00735_),
    .B(_00761_),
    .X(_00762_));
 sky130_fd_sc_hd__nand2_1 _06582_ (.A(net61),
    .B(net13),
    .Y(_00763_));
 sky130_fd_sc_hd__and3_1 _06583_ (.A(net61),
    .B(net13),
    .C(_00762_),
    .X(_00764_));
 sky130_fd_sc_hd__xnor2_1 _06584_ (.A(_00762_),
    .B(_00763_),
    .Y(_00765_));
 sky130_fd_sc_hd__xor2_1 _06585_ (.A(_00734_),
    .B(_00765_),
    .X(_00767_));
 sky130_fd_sc_hd__nand2_1 _06586_ (.A(net62),
    .B(net11),
    .Y(_00768_));
 sky130_fd_sc_hd__and3_1 _06587_ (.A(net62),
    .B(net11),
    .C(_00767_),
    .X(_00769_));
 sky130_fd_sc_hd__xnor2_1 _06588_ (.A(_00767_),
    .B(_00768_),
    .Y(_00770_));
 sky130_fd_sc_hd__xnor2_1 _06589_ (.A(_00732_),
    .B(_00770_),
    .Y(_00771_));
 sky130_fd_sc_hd__nand2_1 _06590_ (.A(net63),
    .B(net10),
    .Y(_00772_));
 sky130_fd_sc_hd__nor2_1 _06591_ (.A(_00771_),
    .B(_00772_),
    .Y(_00773_));
 sky130_fd_sc_hd__xor2_1 _06592_ (.A(_00771_),
    .B(_00772_),
    .X(_00774_));
 sky130_fd_sc_hd__xnor2_1 _06593_ (.A(_00731_),
    .B(_00774_),
    .Y(_00775_));
 sky130_fd_sc_hd__nand2_1 _06594_ (.A(net64),
    .B(net9),
    .Y(_00776_));
 sky130_fd_sc_hd__nor2_1 _06595_ (.A(_00775_),
    .B(_00776_),
    .Y(_00778_));
 sky130_fd_sc_hd__xor2_1 _06596_ (.A(_00775_),
    .B(_00776_),
    .X(_00779_));
 sky130_fd_sc_hd__xnor2_1 _06597_ (.A(_00730_),
    .B(_00779_),
    .Y(_00780_));
 sky130_fd_sc_hd__nand2_1 _06598_ (.A(net34),
    .B(net8),
    .Y(_00781_));
 sky130_fd_sc_hd__nor2_1 _06599_ (.A(_00780_),
    .B(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__xor2_1 _06600_ (.A(_00780_),
    .B(_00781_),
    .X(_00783_));
 sky130_fd_sc_hd__xnor2_1 _06601_ (.A(_00729_),
    .B(_00783_),
    .Y(_00784_));
 sky130_fd_sc_hd__nand2_1 _06602_ (.A(net35),
    .B(net7),
    .Y(_00785_));
 sky130_fd_sc_hd__nor2_1 _06603_ (.A(_00784_),
    .B(_00785_),
    .Y(_00786_));
 sky130_fd_sc_hd__xor2_1 _06604_ (.A(_00784_),
    .B(_00785_),
    .X(_00787_));
 sky130_fd_sc_hd__xnor2_1 _06605_ (.A(_00728_),
    .B(_00787_),
    .Y(_00789_));
 sky130_fd_sc_hd__nand2_1 _06606_ (.A(net36),
    .B(net6),
    .Y(_00790_));
 sky130_fd_sc_hd__nor2_1 _06607_ (.A(_00789_),
    .B(_00790_),
    .Y(_00791_));
 sky130_fd_sc_hd__xor2_1 _06608_ (.A(_00789_),
    .B(_00790_),
    .X(_00792_));
 sky130_fd_sc_hd__xnor2_1 _06609_ (.A(_00727_),
    .B(_00792_),
    .Y(_00793_));
 sky130_fd_sc_hd__nand2_1 _06610_ (.A(net5),
    .B(net37),
    .Y(_00794_));
 sky130_fd_sc_hd__nor2_1 _06611_ (.A(_00793_),
    .B(_00794_),
    .Y(_00795_));
 sky130_fd_sc_hd__xor2_1 _06612_ (.A(_00793_),
    .B(_00794_),
    .X(_00796_));
 sky130_fd_sc_hd__xnor2_1 _06613_ (.A(_00726_),
    .B(_00796_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand2_1 _06614_ (.A(net4),
    .B(net38),
    .Y(_00798_));
 sky130_fd_sc_hd__nor2_1 _06615_ (.A(_00797_),
    .B(_00798_),
    .Y(_00800_));
 sky130_fd_sc_hd__xor2_1 _06616_ (.A(_00797_),
    .B(_00798_),
    .X(_00801_));
 sky130_fd_sc_hd__xnor2_1 _06617_ (.A(_00725_),
    .B(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hd__nand2_1 _06618_ (.A(net3),
    .B(net39),
    .Y(_00803_));
 sky130_fd_sc_hd__nor2_1 _06619_ (.A(_00802_),
    .B(_00803_),
    .Y(_00804_));
 sky130_fd_sc_hd__xor2_1 _06620_ (.A(_00802_),
    .B(_00803_),
    .X(_00805_));
 sky130_fd_sc_hd__xnor2_1 _06621_ (.A(_00724_),
    .B(_00805_),
    .Y(_00806_));
 sky130_fd_sc_hd__nand2_1 _06622_ (.A(net2),
    .B(net40),
    .Y(_00807_));
 sky130_fd_sc_hd__nor2_1 _06623_ (.A(_00806_),
    .B(_00807_),
    .Y(_00808_));
 sky130_fd_sc_hd__xor2_1 _06624_ (.A(_00806_),
    .B(_00807_),
    .X(_00809_));
 sky130_fd_sc_hd__xnor2_1 _06625_ (.A(_00723_),
    .B(_00809_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand2_1 _06626_ (.A(net32),
    .B(net41),
    .Y(_00812_));
 sky130_fd_sc_hd__nor2_1 _06627_ (.A(_00811_),
    .B(_00812_),
    .Y(_00813_));
 sky130_fd_sc_hd__xor2_1 _06628_ (.A(_00811_),
    .B(_00812_),
    .X(_00814_));
 sky130_fd_sc_hd__xnor2_1 _06629_ (.A(_00721_),
    .B(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_1 _06630_ (.A(net31),
    .B(net42),
    .Y(_00816_));
 sky130_fd_sc_hd__nor2_1 _06631_ (.A(_00815_),
    .B(_00816_),
    .Y(_00817_));
 sky130_fd_sc_hd__xor2_1 _06632_ (.A(_00815_),
    .B(_00816_),
    .X(_00818_));
 sky130_fd_sc_hd__xnor2_1 _06633_ (.A(_00720_),
    .B(_00818_),
    .Y(_00819_));
 sky130_fd_sc_hd__nand2_1 _06634_ (.A(net30),
    .B(net43),
    .Y(_00820_));
 sky130_fd_sc_hd__nor2_1 _06635_ (.A(_00819_),
    .B(_00820_),
    .Y(_00822_));
 sky130_fd_sc_hd__xor2_1 _06636_ (.A(_00819_),
    .B(_00820_),
    .X(_00823_));
 sky130_fd_sc_hd__xnor2_1 _06637_ (.A(_00719_),
    .B(_00823_),
    .Y(_00824_));
 sky130_fd_sc_hd__nand2_1 _06638_ (.A(net29),
    .B(net45),
    .Y(_00825_));
 sky130_fd_sc_hd__nor2_1 _06639_ (.A(_00824_),
    .B(_00825_),
    .Y(_00826_));
 sky130_fd_sc_hd__xor2_1 _06640_ (.A(_00824_),
    .B(_00825_),
    .X(_00827_));
 sky130_fd_sc_hd__xnor2_1 _06641_ (.A(_00718_),
    .B(_00827_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand2_1 _06642_ (.A(net28),
    .B(net46),
    .Y(_00829_));
 sky130_fd_sc_hd__nor2_1 _06643_ (.A(_00828_),
    .B(_00829_),
    .Y(_00830_));
 sky130_fd_sc_hd__xor2_1 _06644_ (.A(_00828_),
    .B(_00829_),
    .X(_00831_));
 sky130_fd_sc_hd__xnor2_1 _06645_ (.A(_00717_),
    .B(_00831_),
    .Y(_00833_));
 sky130_fd_sc_hd__nand2_1 _06646_ (.A(net27),
    .B(net47),
    .Y(_00834_));
 sky130_fd_sc_hd__nor2_1 _06647_ (.A(_00833_),
    .B(_00834_),
    .Y(_00835_));
 sky130_fd_sc_hd__xor2_1 _06648_ (.A(_00833_),
    .B(_00834_),
    .X(_00836_));
 sky130_fd_sc_hd__xnor2_1 _06649_ (.A(_00716_),
    .B(_00836_),
    .Y(_00837_));
 sky130_fd_sc_hd__nand2_1 _06650_ (.A(net26),
    .B(net48),
    .Y(_00838_));
 sky130_fd_sc_hd__nor2_1 _06651_ (.A(_00837_),
    .B(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__xor2_1 _06652_ (.A(_00837_),
    .B(_00838_),
    .X(_00840_));
 sky130_fd_sc_hd__xnor2_1 _06653_ (.A(_00715_),
    .B(_00840_),
    .Y(_00841_));
 sky130_fd_sc_hd__nand2_1 _06654_ (.A(net23),
    .B(net49),
    .Y(_00842_));
 sky130_fd_sc_hd__nor2_1 _06655_ (.A(_00841_),
    .B(_00842_),
    .Y(_00844_));
 sky130_fd_sc_hd__xor2_1 _06656_ (.A(_00841_),
    .B(_00842_),
    .X(_00845_));
 sky130_fd_sc_hd__xnor2_1 _06657_ (.A(_00714_),
    .B(_00845_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand2_1 _06658_ (.A(net12),
    .B(net50),
    .Y(_00847_));
 sky130_fd_sc_hd__nor2_1 _06659_ (.A(_00846_),
    .B(_00847_),
    .Y(_00848_));
 sky130_fd_sc_hd__xor2_1 _06660_ (.A(_00846_),
    .B(_00847_),
    .X(_00849_));
 sky130_fd_sc_hd__xor2_1 _06661_ (.A(_00711_),
    .B(_00849_),
    .X(_00850_));
 sky130_fd_sc_hd__and3_1 _06662_ (.A(net1),
    .B(net51),
    .C(_00850_),
    .X(_00851_));
 sky130_fd_sc_hd__a21oi_1 _06663_ (.A1(net1),
    .A2(net51),
    .B1(_00850_),
    .Y(_00852_));
 sky130_fd_sc_hd__nor2_1 _06664_ (.A(_00851_),
    .B(_00852_),
    .Y(\genblk2[25].rca.ripple_adders[26].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _06665_ (.A1(_00711_),
    .A2(_00849_),
    .B1(_00848_),
    .X(_00854_));
 sky130_fd_sc_hd__a21o_1 _06666_ (.A1(_00714_),
    .A2(_00845_),
    .B1(_00844_),
    .X(_00855_));
 sky130_fd_sc_hd__a21o_1 _06667_ (.A1(_00715_),
    .A2(_00840_),
    .B1(_00839_),
    .X(_00856_));
 sky130_fd_sc_hd__a21o_1 _06668_ (.A1(_00716_),
    .A2(_00836_),
    .B1(_00835_),
    .X(_00857_));
 sky130_fd_sc_hd__a21o_1 _06669_ (.A1(_00717_),
    .A2(_00831_),
    .B1(_00830_),
    .X(_00858_));
 sky130_fd_sc_hd__a21o_1 _06670_ (.A1(_00718_),
    .A2(_00827_),
    .B1(_00826_),
    .X(_00859_));
 sky130_fd_sc_hd__a21o_1 _06671_ (.A1(_00719_),
    .A2(_00823_),
    .B1(_00822_),
    .X(_00860_));
 sky130_fd_sc_hd__a21o_1 _06672_ (.A1(_00720_),
    .A2(_00818_),
    .B1(_00817_),
    .X(_00861_));
 sky130_fd_sc_hd__a21o_1 _06673_ (.A1(_00721_),
    .A2(_00814_),
    .B1(_00813_),
    .X(_00862_));
 sky130_fd_sc_hd__a21o_1 _06674_ (.A1(_00723_),
    .A2(_00809_),
    .B1(_00808_),
    .X(_00863_));
 sky130_fd_sc_hd__a21o_1 _06675_ (.A1(_00724_),
    .A2(_00805_),
    .B1(_00804_),
    .X(_00865_));
 sky130_fd_sc_hd__a21o_1 _06676_ (.A1(_00725_),
    .A2(_00801_),
    .B1(_00800_),
    .X(_00866_));
 sky130_fd_sc_hd__a21o_1 _06677_ (.A1(_00726_),
    .A2(_00796_),
    .B1(_00795_),
    .X(_00867_));
 sky130_fd_sc_hd__a21o_1 _06678_ (.A1(_00727_),
    .A2(_00792_),
    .B1(_00791_),
    .X(_00868_));
 sky130_fd_sc_hd__a21o_1 _06679_ (.A1(_00728_),
    .A2(_00787_),
    .B1(_00786_),
    .X(_00869_));
 sky130_fd_sc_hd__a21o_1 _06680_ (.A1(_00729_),
    .A2(_00783_),
    .B1(_00782_),
    .X(_00870_));
 sky130_fd_sc_hd__a21o_1 _06681_ (.A1(_00730_),
    .A2(_00779_),
    .B1(_00778_),
    .X(_00871_));
 sky130_fd_sc_hd__a21o_1 _06682_ (.A1(_00731_),
    .A2(_00774_),
    .B1(_00773_),
    .X(_00872_));
 sky130_fd_sc_hd__a21o_1 _06683_ (.A1(_00732_),
    .A2(_00770_),
    .B1(_00769_),
    .X(_00873_));
 sky130_fd_sc_hd__a21o_1 _06684_ (.A1(_00734_),
    .A2(_00765_),
    .B1(_00764_),
    .X(_00874_));
 sky130_fd_sc_hd__a21o_1 _06685_ (.A1(_00735_),
    .A2(_00761_),
    .B1(_00760_),
    .X(_00876_));
 sky130_fd_sc_hd__a21o_1 _06686_ (.A1(_00736_),
    .A2(_00757_),
    .B1(_00756_),
    .X(_00877_));
 sky130_fd_sc_hd__a21o_1 _06687_ (.A1(_00737_),
    .A2(_00752_),
    .B1(_00751_),
    .X(_00878_));
 sky130_fd_sc_hd__a21o_1 _06688_ (.A1(_00738_),
    .A2(_00747_),
    .B1(_00746_),
    .X(_00879_));
 sky130_fd_sc_hd__a22o_1 _06689_ (.A1(net44),
    .A2(net19),
    .B1(net20),
    .B2(net33),
    .X(_00880_));
 sky130_fd_sc_hd__and3_1 _06690_ (.A(net44),
    .B(net19),
    .C(net20),
    .X(_00881_));
 sky130_fd_sc_hd__a21bo_1 _06691_ (.A1(net33),
    .A2(_00881_),
    .B1_N(_00880_),
    .X(_00882_));
 sky130_fd_sc_hd__a22o_1 _06692_ (.A1(net33),
    .A2(_00740_),
    .B1(_00742_),
    .B2(_00739_),
    .X(_00883_));
 sky130_fd_sc_hd__xnor2_1 _06693_ (.A(_00882_),
    .B(_00883_),
    .Y(_00884_));
 sky130_fd_sc_hd__nand2_1 _06694_ (.A(net55),
    .B(net18),
    .Y(_00885_));
 sky130_fd_sc_hd__and3_1 _06695_ (.A(net55),
    .B(net18),
    .C(_00884_),
    .X(_00887_));
 sky130_fd_sc_hd__nand2b_1 _06696_ (.A_N(_00884_),
    .B(_00885_),
    .Y(_00888_));
 sky130_fd_sc_hd__xor2_1 _06697_ (.A(_00884_),
    .B(_00885_),
    .X(_00889_));
 sky130_fd_sc_hd__xnor2_1 _06698_ (.A(_00879_),
    .B(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__nand2_1 _06699_ (.A(net58),
    .B(net17),
    .Y(_00891_));
 sky130_fd_sc_hd__and3_1 _06700_ (.A(net58),
    .B(net17),
    .C(_00890_),
    .X(_00892_));
 sky130_fd_sc_hd__xnor2_1 _06701_ (.A(_00890_),
    .B(_00891_),
    .Y(_00893_));
 sky130_fd_sc_hd__xor2_1 _06702_ (.A(_00878_),
    .B(_00893_),
    .X(_00894_));
 sky130_fd_sc_hd__nand2_1 _06703_ (.A(net59),
    .B(net16),
    .Y(_00895_));
 sky130_fd_sc_hd__and3_1 _06704_ (.A(net59),
    .B(net16),
    .C(_00894_),
    .X(_00896_));
 sky130_fd_sc_hd__xnor2_1 _06705_ (.A(_00894_),
    .B(_00895_),
    .Y(_00898_));
 sky130_fd_sc_hd__xor2_1 _06706_ (.A(_00877_),
    .B(_00898_),
    .X(_00899_));
 sky130_fd_sc_hd__nand2_1 _06707_ (.A(net60),
    .B(net15),
    .Y(_00900_));
 sky130_fd_sc_hd__and3_1 _06708_ (.A(net60),
    .B(net15),
    .C(_00899_),
    .X(_00901_));
 sky130_fd_sc_hd__xnor2_1 _06709_ (.A(_00899_),
    .B(_00900_),
    .Y(_00902_));
 sky130_fd_sc_hd__xor2_1 _06710_ (.A(_00876_),
    .B(_00902_),
    .X(_00903_));
 sky130_fd_sc_hd__nand2_1 _06711_ (.A(net61),
    .B(net14),
    .Y(_00904_));
 sky130_fd_sc_hd__and3_1 _06712_ (.A(net61),
    .B(net14),
    .C(_00903_),
    .X(_00905_));
 sky130_fd_sc_hd__xnor2_1 _06713_ (.A(_00903_),
    .B(_00904_),
    .Y(_00906_));
 sky130_fd_sc_hd__xor2_1 _06714_ (.A(_00874_),
    .B(_00906_),
    .X(_00907_));
 sky130_fd_sc_hd__nand2_1 _06715_ (.A(net62),
    .B(net13),
    .Y(_00909_));
 sky130_fd_sc_hd__and3_1 _06716_ (.A(net62),
    .B(net13),
    .C(_00907_),
    .X(_00910_));
 sky130_fd_sc_hd__xnor2_1 _06717_ (.A(_00907_),
    .B(_00909_),
    .Y(_00911_));
 sky130_fd_sc_hd__xnor2_1 _06718_ (.A(_00873_),
    .B(_00911_),
    .Y(_00912_));
 sky130_fd_sc_hd__nand2_1 _06719_ (.A(net63),
    .B(net11),
    .Y(_00913_));
 sky130_fd_sc_hd__nor2_1 _06720_ (.A(_00912_),
    .B(_00913_),
    .Y(_00914_));
 sky130_fd_sc_hd__xor2_1 _06721_ (.A(_00912_),
    .B(_00913_),
    .X(_00915_));
 sky130_fd_sc_hd__xnor2_1 _06722_ (.A(_00872_),
    .B(_00915_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand2_1 _06723_ (.A(net64),
    .B(net10),
    .Y(_00917_));
 sky130_fd_sc_hd__nor2_1 _06724_ (.A(_00916_),
    .B(_00917_),
    .Y(_00918_));
 sky130_fd_sc_hd__xor2_1 _06725_ (.A(_00916_),
    .B(_00917_),
    .X(_00920_));
 sky130_fd_sc_hd__xnor2_1 _06726_ (.A(_00871_),
    .B(_00920_),
    .Y(_00921_));
 sky130_fd_sc_hd__nand2_1 _06727_ (.A(net34),
    .B(net9),
    .Y(_00922_));
 sky130_fd_sc_hd__nor2_1 _06728_ (.A(_00921_),
    .B(_00922_),
    .Y(_00923_));
 sky130_fd_sc_hd__xor2_1 _06729_ (.A(_00921_),
    .B(_00922_),
    .X(_00924_));
 sky130_fd_sc_hd__xnor2_1 _06730_ (.A(_00870_),
    .B(_00924_),
    .Y(_00925_));
 sky130_fd_sc_hd__nand2_1 _06731_ (.A(net35),
    .B(net8),
    .Y(_00926_));
 sky130_fd_sc_hd__nor2_1 _06732_ (.A(_00925_),
    .B(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hd__xor2_1 _06733_ (.A(_00925_),
    .B(_00926_),
    .X(_00928_));
 sky130_fd_sc_hd__xnor2_1 _06734_ (.A(_00869_),
    .B(_00928_),
    .Y(_00929_));
 sky130_fd_sc_hd__nand2_1 _06735_ (.A(net36),
    .B(net7),
    .Y(_00931_));
 sky130_fd_sc_hd__nor2_1 _06736_ (.A(_00929_),
    .B(_00931_),
    .Y(_00932_));
 sky130_fd_sc_hd__xor2_1 _06737_ (.A(_00929_),
    .B(_00931_),
    .X(_00933_));
 sky130_fd_sc_hd__xnor2_1 _06738_ (.A(_00868_),
    .B(_00933_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand2_1 _06739_ (.A(net37),
    .B(net6),
    .Y(_00935_));
 sky130_fd_sc_hd__nor2_1 _06740_ (.A(_00934_),
    .B(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__xor2_1 _06741_ (.A(_00934_),
    .B(_00935_),
    .X(_00937_));
 sky130_fd_sc_hd__xnor2_1 _06742_ (.A(_00867_),
    .B(_00937_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_1 _06743_ (.A(net5),
    .B(net38),
    .Y(_00939_));
 sky130_fd_sc_hd__nor2_1 _06744_ (.A(_00938_),
    .B(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__xor2_1 _06745_ (.A(_00938_),
    .B(_00939_),
    .X(_00942_));
 sky130_fd_sc_hd__xnor2_1 _06746_ (.A(_00866_),
    .B(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__nand2_1 _06747_ (.A(net4),
    .B(net39),
    .Y(_00944_));
 sky130_fd_sc_hd__nor2_1 _06748_ (.A(_00943_),
    .B(_00944_),
    .Y(_00945_));
 sky130_fd_sc_hd__xor2_1 _06749_ (.A(_00943_),
    .B(_00944_),
    .X(_00946_));
 sky130_fd_sc_hd__xnor2_1 _06750_ (.A(_00865_),
    .B(_00946_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand2_1 _06751_ (.A(net3),
    .B(net40),
    .Y(_00948_));
 sky130_fd_sc_hd__nor2_1 _06752_ (.A(_00947_),
    .B(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__xor2_1 _06753_ (.A(_00947_),
    .B(_00948_),
    .X(_00950_));
 sky130_fd_sc_hd__xnor2_1 _06754_ (.A(_00863_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__nand2_1 _06755_ (.A(net2),
    .B(net41),
    .Y(_00953_));
 sky130_fd_sc_hd__nor2_1 _06756_ (.A(_00951_),
    .B(_00953_),
    .Y(_00954_));
 sky130_fd_sc_hd__xor2_1 _06757_ (.A(_00951_),
    .B(_00953_),
    .X(_00955_));
 sky130_fd_sc_hd__xnor2_1 _06758_ (.A(_00862_),
    .B(_00955_),
    .Y(_00956_));
 sky130_fd_sc_hd__nand2_1 _06759_ (.A(net32),
    .B(net42),
    .Y(_00957_));
 sky130_fd_sc_hd__nor2_1 _06760_ (.A(_00956_),
    .B(_00957_),
    .Y(_00958_));
 sky130_fd_sc_hd__xor2_1 _06761_ (.A(_00956_),
    .B(_00957_),
    .X(_00959_));
 sky130_fd_sc_hd__xnor2_1 _06762_ (.A(_00861_),
    .B(_00959_),
    .Y(_00960_));
 sky130_fd_sc_hd__nand2_1 _06763_ (.A(net31),
    .B(net43),
    .Y(_00961_));
 sky130_fd_sc_hd__nor2_1 _06764_ (.A(_00960_),
    .B(_00961_),
    .Y(_00962_));
 sky130_fd_sc_hd__xor2_1 _06765_ (.A(_00960_),
    .B(_00961_),
    .X(_00964_));
 sky130_fd_sc_hd__xnor2_1 _06766_ (.A(_00860_),
    .B(_00964_),
    .Y(_00965_));
 sky130_fd_sc_hd__nand2_1 _06767_ (.A(net30),
    .B(net45),
    .Y(_00966_));
 sky130_fd_sc_hd__nor2_1 _06768_ (.A(_00965_),
    .B(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__xor2_1 _06769_ (.A(_00965_),
    .B(_00966_),
    .X(_00968_));
 sky130_fd_sc_hd__xnor2_1 _06770_ (.A(_00859_),
    .B(_00968_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_1 _06771_ (.A(net29),
    .B(net46),
    .Y(_00970_));
 sky130_fd_sc_hd__nor2_1 _06772_ (.A(_00969_),
    .B(_00970_),
    .Y(_00971_));
 sky130_fd_sc_hd__xor2_1 _06773_ (.A(_00969_),
    .B(_00970_),
    .X(_00972_));
 sky130_fd_sc_hd__xnor2_1 _06774_ (.A(_00858_),
    .B(_00972_),
    .Y(_00973_));
 sky130_fd_sc_hd__nand2_1 _06775_ (.A(net28),
    .B(net47),
    .Y(_00975_));
 sky130_fd_sc_hd__nor2_1 _06776_ (.A(_00973_),
    .B(_00975_),
    .Y(_00976_));
 sky130_fd_sc_hd__xor2_1 _06777_ (.A(_00973_),
    .B(_00975_),
    .X(_00977_));
 sky130_fd_sc_hd__xnor2_1 _06778_ (.A(_00857_),
    .B(_00977_),
    .Y(_00978_));
 sky130_fd_sc_hd__nand2_1 _06779_ (.A(net27),
    .B(net48),
    .Y(_00979_));
 sky130_fd_sc_hd__nor2_1 _06780_ (.A(_00978_),
    .B(_00979_),
    .Y(_00980_));
 sky130_fd_sc_hd__xor2_1 _06781_ (.A(_00978_),
    .B(_00979_),
    .X(_00981_));
 sky130_fd_sc_hd__xnor2_1 _06782_ (.A(_00856_),
    .B(_00981_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2_1 _06783_ (.A(net26),
    .B(net49),
    .Y(_00983_));
 sky130_fd_sc_hd__nor2_1 _06784_ (.A(_00982_),
    .B(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__xor2_1 _06785_ (.A(_00982_),
    .B(_00983_),
    .X(_00986_));
 sky130_fd_sc_hd__xnor2_1 _06786_ (.A(_00855_),
    .B(_00986_),
    .Y(_00987_));
 sky130_fd_sc_hd__nand2_1 _06787_ (.A(net23),
    .B(net50),
    .Y(_00988_));
 sky130_fd_sc_hd__nor2_1 _06788_ (.A(_00987_),
    .B(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__xor2_1 _06789_ (.A(_00987_),
    .B(_00988_),
    .X(_00990_));
 sky130_fd_sc_hd__xnor2_1 _06790_ (.A(_00854_),
    .B(_00990_),
    .Y(_00991_));
 sky130_fd_sc_hd__nand2_1 _06791_ (.A(net12),
    .B(net51),
    .Y(_00992_));
 sky130_fd_sc_hd__nor2_1 _06792_ (.A(_00991_),
    .B(_00992_),
    .Y(_00993_));
 sky130_fd_sc_hd__xor2_1 _06793_ (.A(_00991_),
    .B(_00992_),
    .X(_00994_));
 sky130_fd_sc_hd__xor2_1 _06794_ (.A(_00851_),
    .B(_00994_),
    .X(_00995_));
 sky130_fd_sc_hd__and3_1 _06795_ (.A(net1),
    .B(net52),
    .C(_00995_),
    .X(_00997_));
 sky130_fd_sc_hd__a21oi_1 _06796_ (.A1(net1),
    .A2(net52),
    .B1(_00995_),
    .Y(_00998_));
 sky130_fd_sc_hd__nor2_1 _06797_ (.A(_00997_),
    .B(_00998_),
    .Y(\genblk2[26].rca.ripple_adders[27].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _06798_ (.A1(_00851_),
    .A2(_00994_),
    .B1(_00993_),
    .X(_00999_));
 sky130_fd_sc_hd__a21o_1 _06799_ (.A1(_00854_),
    .A2(_00990_),
    .B1(_00989_),
    .X(_01000_));
 sky130_fd_sc_hd__a21o_1 _06800_ (.A1(_00855_),
    .A2(_00986_),
    .B1(_00984_),
    .X(_01001_));
 sky130_fd_sc_hd__a21o_1 _06801_ (.A1(_00856_),
    .A2(_00981_),
    .B1(_00980_),
    .X(_01002_));
 sky130_fd_sc_hd__a21o_1 _06802_ (.A1(_00857_),
    .A2(_00977_),
    .B1(_00976_),
    .X(_01003_));
 sky130_fd_sc_hd__a21o_1 _06803_ (.A1(_00858_),
    .A2(_00972_),
    .B1(_00971_),
    .X(_01004_));
 sky130_fd_sc_hd__a21o_1 _06804_ (.A1(_00859_),
    .A2(_00968_),
    .B1(_00967_),
    .X(_01005_));
 sky130_fd_sc_hd__a21o_1 _06805_ (.A1(_00860_),
    .A2(_00964_),
    .B1(_00962_),
    .X(_01007_));
 sky130_fd_sc_hd__a21o_1 _06806_ (.A1(_00861_),
    .A2(_00959_),
    .B1(_00958_),
    .X(_01008_));
 sky130_fd_sc_hd__a21o_1 _06807_ (.A1(_00862_),
    .A2(_00955_),
    .B1(_00954_),
    .X(_01009_));
 sky130_fd_sc_hd__a21o_1 _06808_ (.A1(_00863_),
    .A2(_00950_),
    .B1(_00949_),
    .X(_01010_));
 sky130_fd_sc_hd__a21o_1 _06809_ (.A1(_00865_),
    .A2(_00946_),
    .B1(_00945_),
    .X(_01011_));
 sky130_fd_sc_hd__a21o_1 _06810_ (.A1(_00866_),
    .A2(_00942_),
    .B1(_00940_),
    .X(_01012_));
 sky130_fd_sc_hd__a21o_1 _06811_ (.A1(_00867_),
    .A2(_00937_),
    .B1(_00936_),
    .X(_01013_));
 sky130_fd_sc_hd__a21o_1 _06812_ (.A1(_00868_),
    .A2(_00933_),
    .B1(_00932_),
    .X(_01014_));
 sky130_fd_sc_hd__a21o_1 _06813_ (.A1(_00869_),
    .A2(_00928_),
    .B1(_00927_),
    .X(_01015_));
 sky130_fd_sc_hd__a21o_1 _06814_ (.A1(_00870_),
    .A2(_00924_),
    .B1(_00923_),
    .X(_01016_));
 sky130_fd_sc_hd__a21o_1 _06815_ (.A1(_00871_),
    .A2(_00920_),
    .B1(_00918_),
    .X(_01018_));
 sky130_fd_sc_hd__a21o_1 _06816_ (.A1(_00872_),
    .A2(_00915_),
    .B1(_00914_),
    .X(_01019_));
 sky130_fd_sc_hd__a21o_1 _06817_ (.A1(_00873_),
    .A2(_00911_),
    .B1(_00910_),
    .X(_01020_));
 sky130_fd_sc_hd__a21o_1 _06818_ (.A1(_00874_),
    .A2(_00906_),
    .B1(_00905_),
    .X(_01021_));
 sky130_fd_sc_hd__a21o_1 _06819_ (.A1(_00876_),
    .A2(_00902_),
    .B1(_00901_),
    .X(_01022_));
 sky130_fd_sc_hd__a21o_1 _06820_ (.A1(_00877_),
    .A2(_00898_),
    .B1(_00896_),
    .X(_01023_));
 sky130_fd_sc_hd__a21o_1 _06821_ (.A1(_00878_),
    .A2(_00893_),
    .B1(_00892_),
    .X(_01024_));
 sky130_fd_sc_hd__a21o_1 _06822_ (.A1(_00879_),
    .A2(_00888_),
    .B1(_00887_),
    .X(_01025_));
 sky130_fd_sc_hd__a22o_1 _06823_ (.A1(net44),
    .A2(net20),
    .B1(net21),
    .B2(net33),
    .X(_01026_));
 sky130_fd_sc_hd__and3_1 _06824_ (.A(net44),
    .B(net20),
    .C(net21),
    .X(_01027_));
 sky130_fd_sc_hd__a21bo_1 _06825_ (.A1(net33),
    .A2(_01027_),
    .B1_N(_01026_),
    .X(_01029_));
 sky130_fd_sc_hd__a22o_1 _06826_ (.A1(net33),
    .A2(_00881_),
    .B1(_00883_),
    .B2(_00880_),
    .X(_01030_));
 sky130_fd_sc_hd__xnor2_1 _06827_ (.A(_01029_),
    .B(_01030_),
    .Y(_01031_));
 sky130_fd_sc_hd__nand2_1 _06828_ (.A(net55),
    .B(net19),
    .Y(_01032_));
 sky130_fd_sc_hd__and3_1 _06829_ (.A(net55),
    .B(net19),
    .C(_01031_),
    .X(_01033_));
 sky130_fd_sc_hd__nand2b_1 _06830_ (.A_N(_01031_),
    .B(_01032_),
    .Y(_01034_));
 sky130_fd_sc_hd__xor2_1 _06831_ (.A(_01031_),
    .B(_01032_),
    .X(_01035_));
 sky130_fd_sc_hd__xnor2_1 _06832_ (.A(_01025_),
    .B(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hd__nand2_1 _06833_ (.A(net58),
    .B(net18),
    .Y(_01037_));
 sky130_fd_sc_hd__and3_1 _06834_ (.A(net58),
    .B(net18),
    .C(_01036_),
    .X(_01038_));
 sky130_fd_sc_hd__xnor2_1 _06835_ (.A(_01036_),
    .B(_01037_),
    .Y(_01040_));
 sky130_fd_sc_hd__xor2_1 _06836_ (.A(_01024_),
    .B(_01040_),
    .X(_01041_));
 sky130_fd_sc_hd__nand2_1 _06837_ (.A(net59),
    .B(net17),
    .Y(_01042_));
 sky130_fd_sc_hd__and3_1 _06838_ (.A(net59),
    .B(net17),
    .C(_01041_),
    .X(_01043_));
 sky130_fd_sc_hd__xnor2_1 _06839_ (.A(_01041_),
    .B(_01042_),
    .Y(_01044_));
 sky130_fd_sc_hd__xor2_1 _06840_ (.A(_01023_),
    .B(_01044_),
    .X(_01045_));
 sky130_fd_sc_hd__nand2_1 _06841_ (.A(net60),
    .B(net16),
    .Y(_01046_));
 sky130_fd_sc_hd__and3_1 _06842_ (.A(net60),
    .B(net16),
    .C(_01045_),
    .X(_01047_));
 sky130_fd_sc_hd__xnor2_1 _06843_ (.A(_01045_),
    .B(_01046_),
    .Y(_01048_));
 sky130_fd_sc_hd__xor2_1 _06844_ (.A(_01022_),
    .B(_01048_),
    .X(_01049_));
 sky130_fd_sc_hd__nand2_1 _06845_ (.A(net61),
    .B(net15),
    .Y(_01051_));
 sky130_fd_sc_hd__and3_1 _06846_ (.A(net61),
    .B(net15),
    .C(_01049_),
    .X(_01052_));
 sky130_fd_sc_hd__xnor2_1 _06847_ (.A(_01049_),
    .B(_01051_),
    .Y(_01053_));
 sky130_fd_sc_hd__xnor2_1 _06848_ (.A(_01021_),
    .B(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__nand2_1 _06849_ (.A(net62),
    .B(net14),
    .Y(_01055_));
 sky130_fd_sc_hd__nor2_1 _06850_ (.A(_01054_),
    .B(_01055_),
    .Y(_01056_));
 sky130_fd_sc_hd__xor2_1 _06851_ (.A(_01054_),
    .B(_01055_),
    .X(_01057_));
 sky130_fd_sc_hd__xnor2_1 _06852_ (.A(_01020_),
    .B(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__nand2_1 _06853_ (.A(net63),
    .B(net13),
    .Y(_01059_));
 sky130_fd_sc_hd__nor2_1 _06854_ (.A(_01058_),
    .B(_01059_),
    .Y(_01060_));
 sky130_fd_sc_hd__xor2_1 _06855_ (.A(_01058_),
    .B(_01059_),
    .X(_01062_));
 sky130_fd_sc_hd__xnor2_1 _06856_ (.A(_01019_),
    .B(_01062_),
    .Y(_01063_));
 sky130_fd_sc_hd__nand2_1 _06857_ (.A(net64),
    .B(net11),
    .Y(_01064_));
 sky130_fd_sc_hd__nor2_1 _06858_ (.A(_01063_),
    .B(_01064_),
    .Y(_01065_));
 sky130_fd_sc_hd__xor2_1 _06859_ (.A(_01063_),
    .B(_01064_),
    .X(_01066_));
 sky130_fd_sc_hd__xnor2_1 _06860_ (.A(_01018_),
    .B(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand2_1 _06861_ (.A(net34),
    .B(net10),
    .Y(_01068_));
 sky130_fd_sc_hd__nor2_1 _06862_ (.A(_01067_),
    .B(_01068_),
    .Y(_01069_));
 sky130_fd_sc_hd__xor2_1 _06863_ (.A(_01067_),
    .B(_01068_),
    .X(_01070_));
 sky130_fd_sc_hd__xnor2_1 _06864_ (.A(_01016_),
    .B(_01070_),
    .Y(_01071_));
 sky130_fd_sc_hd__nand2_1 _06865_ (.A(net35),
    .B(net9),
    .Y(_01073_));
 sky130_fd_sc_hd__nor2_1 _06866_ (.A(_01071_),
    .B(_01073_),
    .Y(_01074_));
 sky130_fd_sc_hd__xor2_1 _06867_ (.A(_01071_),
    .B(_01073_),
    .X(_01075_));
 sky130_fd_sc_hd__xnor2_1 _06868_ (.A(_01015_),
    .B(_01075_),
    .Y(_01076_));
 sky130_fd_sc_hd__nand2_1 _06869_ (.A(net36),
    .B(net8),
    .Y(_01077_));
 sky130_fd_sc_hd__nor2_1 _06870_ (.A(_01076_),
    .B(_01077_),
    .Y(_01078_));
 sky130_fd_sc_hd__xor2_1 _06871_ (.A(_01076_),
    .B(_01077_),
    .X(_01079_));
 sky130_fd_sc_hd__xnor2_1 _06872_ (.A(_01014_),
    .B(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__nand2_1 _06873_ (.A(net37),
    .B(net7),
    .Y(_01081_));
 sky130_fd_sc_hd__nor2_1 _06874_ (.A(_01080_),
    .B(_01081_),
    .Y(_01082_));
 sky130_fd_sc_hd__xor2_1 _06875_ (.A(_01080_),
    .B(_01081_),
    .X(_01084_));
 sky130_fd_sc_hd__xnor2_1 _06876_ (.A(_01013_),
    .B(_01084_),
    .Y(_01085_));
 sky130_fd_sc_hd__nand2_1 _06877_ (.A(net6),
    .B(net38),
    .Y(_01086_));
 sky130_fd_sc_hd__nor2_1 _06878_ (.A(_01085_),
    .B(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hd__xor2_1 _06879_ (.A(_01085_),
    .B(_01086_),
    .X(_01088_));
 sky130_fd_sc_hd__xnor2_1 _06880_ (.A(_01012_),
    .B(_01088_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand2_1 _06881_ (.A(net5),
    .B(net39),
    .Y(_01090_));
 sky130_fd_sc_hd__nor2_1 _06882_ (.A(_01089_),
    .B(_01090_),
    .Y(_01091_));
 sky130_fd_sc_hd__xor2_1 _06883_ (.A(_01089_),
    .B(_01090_),
    .X(_01092_));
 sky130_fd_sc_hd__xnor2_1 _06884_ (.A(_01011_),
    .B(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__nand2_1 _06885_ (.A(net4),
    .B(net40),
    .Y(_01095_));
 sky130_fd_sc_hd__nor2_1 _06886_ (.A(_01093_),
    .B(_01095_),
    .Y(_01096_));
 sky130_fd_sc_hd__xor2_1 _06887_ (.A(_01093_),
    .B(_01095_),
    .X(_01097_));
 sky130_fd_sc_hd__xnor2_1 _06888_ (.A(_01010_),
    .B(_01097_),
    .Y(_01098_));
 sky130_fd_sc_hd__nand2_1 _06889_ (.A(net3),
    .B(net41),
    .Y(_01099_));
 sky130_fd_sc_hd__nor2_1 _06890_ (.A(_01098_),
    .B(_01099_),
    .Y(_01100_));
 sky130_fd_sc_hd__xor2_1 _06891_ (.A(_01098_),
    .B(_01099_),
    .X(_01101_));
 sky130_fd_sc_hd__xnor2_1 _06892_ (.A(_01009_),
    .B(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__nand2_1 _06893_ (.A(net2),
    .B(net42),
    .Y(_01103_));
 sky130_fd_sc_hd__nor2_1 _06894_ (.A(_01102_),
    .B(_01103_),
    .Y(_01104_));
 sky130_fd_sc_hd__xor2_1 _06895_ (.A(_01102_),
    .B(_01103_),
    .X(_01106_));
 sky130_fd_sc_hd__xnor2_1 _06896_ (.A(_01008_),
    .B(_01106_),
    .Y(_01107_));
 sky130_fd_sc_hd__nand2_1 _06897_ (.A(net32),
    .B(net43),
    .Y(_01108_));
 sky130_fd_sc_hd__nor2_1 _06898_ (.A(_01107_),
    .B(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__xor2_1 _06899_ (.A(_01107_),
    .B(_01108_),
    .X(_01110_));
 sky130_fd_sc_hd__xnor2_1 _06900_ (.A(_01007_),
    .B(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__nand2_1 _06901_ (.A(net31),
    .B(net45),
    .Y(_01112_));
 sky130_fd_sc_hd__nor2_1 _06902_ (.A(_01111_),
    .B(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__xor2_1 _06903_ (.A(_01111_),
    .B(_01112_),
    .X(_01114_));
 sky130_fd_sc_hd__xnor2_1 _06904_ (.A(_01005_),
    .B(_01114_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand2_1 _06905_ (.A(net30),
    .B(net46),
    .Y(_01117_));
 sky130_fd_sc_hd__nor2_1 _06906_ (.A(_01115_),
    .B(_01117_),
    .Y(_01118_));
 sky130_fd_sc_hd__xor2_1 _06907_ (.A(_01115_),
    .B(_01117_),
    .X(_01119_));
 sky130_fd_sc_hd__xnor2_1 _06908_ (.A(_01004_),
    .B(_01119_),
    .Y(_01120_));
 sky130_fd_sc_hd__nand2_1 _06909_ (.A(net29),
    .B(net47),
    .Y(_01121_));
 sky130_fd_sc_hd__nor2_1 _06910_ (.A(_01120_),
    .B(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__xor2_1 _06911_ (.A(_01120_),
    .B(_01121_),
    .X(_01123_));
 sky130_fd_sc_hd__xnor2_1 _06912_ (.A(_01003_),
    .B(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2_1 _06913_ (.A(net28),
    .B(net48),
    .Y(_01125_));
 sky130_fd_sc_hd__nor2_1 _06914_ (.A(_01124_),
    .B(_01125_),
    .Y(_01126_));
 sky130_fd_sc_hd__xor2_1 _06915_ (.A(_01124_),
    .B(_01125_),
    .X(_01128_));
 sky130_fd_sc_hd__xnor2_1 _06916_ (.A(_01002_),
    .B(_01128_),
    .Y(_01129_));
 sky130_fd_sc_hd__nand2_1 _06917_ (.A(net27),
    .B(net49),
    .Y(_01130_));
 sky130_fd_sc_hd__nor2_1 _06918_ (.A(_01129_),
    .B(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__xor2_1 _06919_ (.A(_01129_),
    .B(_01130_),
    .X(_01132_));
 sky130_fd_sc_hd__xnor2_1 _06920_ (.A(_01001_),
    .B(_01132_),
    .Y(_01133_));
 sky130_fd_sc_hd__nand2_1 _06921_ (.A(net26),
    .B(net50),
    .Y(_01134_));
 sky130_fd_sc_hd__nor2_1 _06922_ (.A(_01133_),
    .B(_01134_),
    .Y(_01135_));
 sky130_fd_sc_hd__xor2_1 _06923_ (.A(_01133_),
    .B(_01134_),
    .X(_01136_));
 sky130_fd_sc_hd__xnor2_1 _06924_ (.A(_01000_),
    .B(_01136_),
    .Y(_01137_));
 sky130_fd_sc_hd__nand2_1 _06925_ (.A(net23),
    .B(net51),
    .Y(_01139_));
 sky130_fd_sc_hd__nor2_1 _06926_ (.A(_01137_),
    .B(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__xor2_1 _06927_ (.A(_01137_),
    .B(_01139_),
    .X(_01141_));
 sky130_fd_sc_hd__xnor2_1 _06928_ (.A(_00999_),
    .B(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__nand2_1 _06929_ (.A(net12),
    .B(net52),
    .Y(_01143_));
 sky130_fd_sc_hd__nor2_1 _06930_ (.A(_01142_),
    .B(_01143_),
    .Y(_01144_));
 sky130_fd_sc_hd__xor2_1 _06931_ (.A(_01142_),
    .B(_01143_),
    .X(_01145_));
 sky130_fd_sc_hd__xor2_1 _06932_ (.A(_00997_),
    .B(_01145_),
    .X(_01146_));
 sky130_fd_sc_hd__and3_1 _06933_ (.A(net1),
    .B(net53),
    .C(_01146_),
    .X(_01147_));
 sky130_fd_sc_hd__a21oi_1 _06934_ (.A1(net1),
    .A2(net53),
    .B1(_01146_),
    .Y(_01148_));
 sky130_fd_sc_hd__nor2_1 _06935_ (.A(_01147_),
    .B(_01148_),
    .Y(\genblk2[27].rca.ripple_adders[28].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _06936_ (.A1(_00997_),
    .A2(_01145_),
    .B1(_01144_),
    .X(_01150_));
 sky130_fd_sc_hd__a21o_1 _06937_ (.A1(_00999_),
    .A2(_01141_),
    .B1(_01140_),
    .X(_01151_));
 sky130_fd_sc_hd__a21o_1 _06938_ (.A1(_01000_),
    .A2(_01136_),
    .B1(_01135_),
    .X(_01152_));
 sky130_fd_sc_hd__a21o_1 _06939_ (.A1(_01001_),
    .A2(_01132_),
    .B1(_01131_),
    .X(_01153_));
 sky130_fd_sc_hd__a21o_1 _06940_ (.A1(_01002_),
    .A2(_01128_),
    .B1(_01126_),
    .X(_01154_));
 sky130_fd_sc_hd__a21o_1 _06941_ (.A1(_01003_),
    .A2(_01123_),
    .B1(_01122_),
    .X(_01155_));
 sky130_fd_sc_hd__a21o_1 _06942_ (.A1(_01004_),
    .A2(_01119_),
    .B1(_01118_),
    .X(_01156_));
 sky130_fd_sc_hd__a21o_1 _06943_ (.A1(_01005_),
    .A2(_01114_),
    .B1(_01113_),
    .X(_01157_));
 sky130_fd_sc_hd__a21o_1 _06944_ (.A1(_01007_),
    .A2(_01110_),
    .B1(_01109_),
    .X(_01158_));
 sky130_fd_sc_hd__a21o_1 _06945_ (.A1(_01008_),
    .A2(_01106_),
    .B1(_01104_),
    .X(_01160_));
 sky130_fd_sc_hd__a21o_1 _06946_ (.A1(_01009_),
    .A2(_01101_),
    .B1(_01100_),
    .X(_01161_));
 sky130_fd_sc_hd__a21o_1 _06947_ (.A1(_01010_),
    .A2(_01097_),
    .B1(_01096_),
    .X(_01162_));
 sky130_fd_sc_hd__a21o_1 _06948_ (.A1(_01011_),
    .A2(_01092_),
    .B1(_01091_),
    .X(_01163_));
 sky130_fd_sc_hd__a21o_1 _06949_ (.A1(_01012_),
    .A2(_01088_),
    .B1(_01087_),
    .X(_01164_));
 sky130_fd_sc_hd__a21o_1 _06950_ (.A1(_01013_),
    .A2(_01084_),
    .B1(_01082_),
    .X(_01165_));
 sky130_fd_sc_hd__a21o_1 _06951_ (.A1(_01014_),
    .A2(_01079_),
    .B1(_01078_),
    .X(_01166_));
 sky130_fd_sc_hd__a21o_1 _06952_ (.A1(_01015_),
    .A2(_01075_),
    .B1(_01074_),
    .X(_01167_));
 sky130_fd_sc_hd__a21o_1 _06953_ (.A1(_01016_),
    .A2(_01070_),
    .B1(_01069_),
    .X(_01168_));
 sky130_fd_sc_hd__a21o_1 _06954_ (.A1(_01018_),
    .A2(_01066_),
    .B1(_01065_),
    .X(_01169_));
 sky130_fd_sc_hd__a21o_1 _06955_ (.A1(_01019_),
    .A2(_01062_),
    .B1(_01060_),
    .X(_01171_));
 sky130_fd_sc_hd__a21o_1 _06956_ (.A1(_01020_),
    .A2(_01057_),
    .B1(_01056_),
    .X(_01172_));
 sky130_fd_sc_hd__a21o_1 _06957_ (.A1(_01021_),
    .A2(_01053_),
    .B1(_01052_),
    .X(_01173_));
 sky130_fd_sc_hd__a21o_1 _06958_ (.A1(_01022_),
    .A2(_01048_),
    .B1(_01047_),
    .X(_01174_));
 sky130_fd_sc_hd__a21o_1 _06959_ (.A1(_01023_),
    .A2(_01044_),
    .B1(_01043_),
    .X(_01175_));
 sky130_fd_sc_hd__a21o_1 _06960_ (.A1(_01024_),
    .A2(_01040_),
    .B1(_01038_),
    .X(_01176_));
 sky130_fd_sc_hd__a21o_1 _06961_ (.A1(_01025_),
    .A2(_01034_),
    .B1(_01033_),
    .X(_01177_));
 sky130_fd_sc_hd__a22o_1 _06962_ (.A1(net44),
    .A2(net21),
    .B1(net22),
    .B2(net33),
    .X(_01178_));
 sky130_fd_sc_hd__and4_1 _06963_ (.A(net33),
    .B(net44),
    .C(net21),
    .D(net22),
    .X(_01179_));
 sky130_fd_sc_hd__inv_2 _06964_ (.A(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__nand2_1 _06965_ (.A(_01178_),
    .B(_01180_),
    .Y(_01182_));
 sky130_fd_sc_hd__a22o_1 _06966_ (.A1(net33),
    .A2(_01027_),
    .B1(_01030_),
    .B2(_01026_),
    .X(_01183_));
 sky130_fd_sc_hd__xnor2_1 _06967_ (.A(_01182_),
    .B(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__nand2_1 _06968_ (.A(net55),
    .B(net20),
    .Y(_01185_));
 sky130_fd_sc_hd__and3_1 _06969_ (.A(net55),
    .B(net20),
    .C(_01184_),
    .X(_01186_));
 sky130_fd_sc_hd__nand2b_1 _06970_ (.A_N(_01184_),
    .B(_01185_),
    .Y(_01187_));
 sky130_fd_sc_hd__xor2_1 _06971_ (.A(_01184_),
    .B(_01185_),
    .X(_01188_));
 sky130_fd_sc_hd__xnor2_1 _06972_ (.A(_01177_),
    .B(_01188_),
    .Y(_01189_));
 sky130_fd_sc_hd__nand2_1 _06973_ (.A(net58),
    .B(net19),
    .Y(_01190_));
 sky130_fd_sc_hd__and3_1 _06974_ (.A(net58),
    .B(net19),
    .C(_01189_),
    .X(_01191_));
 sky130_fd_sc_hd__xnor2_1 _06975_ (.A(_01189_),
    .B(_01190_),
    .Y(_01193_));
 sky130_fd_sc_hd__xor2_1 _06976_ (.A(_01176_),
    .B(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__nand2_1 _06977_ (.A(net59),
    .B(net18),
    .Y(_01195_));
 sky130_fd_sc_hd__and3_1 _06978_ (.A(net59),
    .B(net18),
    .C(_01194_),
    .X(_01196_));
 sky130_fd_sc_hd__xnor2_1 _06979_ (.A(_01194_),
    .B(_01195_),
    .Y(_01197_));
 sky130_fd_sc_hd__xor2_1 _06980_ (.A(_01175_),
    .B(_01197_),
    .X(_01198_));
 sky130_fd_sc_hd__nand2_1 _06981_ (.A(net60),
    .B(net17),
    .Y(_01199_));
 sky130_fd_sc_hd__and3_1 _06982_ (.A(net60),
    .B(net17),
    .C(_01198_),
    .X(_01200_));
 sky130_fd_sc_hd__xnor2_1 _06983_ (.A(_01198_),
    .B(_01199_),
    .Y(_01201_));
 sky130_fd_sc_hd__xor2_1 _06984_ (.A(_01174_),
    .B(_01201_),
    .X(_01202_));
 sky130_fd_sc_hd__nand2_1 _06985_ (.A(net61),
    .B(net16),
    .Y(_01204_));
 sky130_fd_sc_hd__and3_1 _06986_ (.A(net61),
    .B(net16),
    .C(_01202_),
    .X(_01205_));
 sky130_fd_sc_hd__xnor2_1 _06987_ (.A(_01202_),
    .B(_01204_),
    .Y(_01206_));
 sky130_fd_sc_hd__xnor2_1 _06988_ (.A(_01173_),
    .B(_01206_),
    .Y(_01207_));
 sky130_fd_sc_hd__nand2_1 _06989_ (.A(net62),
    .B(net15),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _06990_ (.A(_01207_),
    .B(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__xor2_1 _06991_ (.A(_01207_),
    .B(_01208_),
    .X(_01210_));
 sky130_fd_sc_hd__xnor2_1 _06992_ (.A(_01172_),
    .B(_01210_),
    .Y(_01211_));
 sky130_fd_sc_hd__nand2_1 _06993_ (.A(net63),
    .B(net14),
    .Y(_01212_));
 sky130_fd_sc_hd__nor2_1 _06994_ (.A(_01211_),
    .B(_01212_),
    .Y(_01213_));
 sky130_fd_sc_hd__xor2_1 _06995_ (.A(_01211_),
    .B(_01212_),
    .X(_01215_));
 sky130_fd_sc_hd__xnor2_1 _06996_ (.A(_01171_),
    .B(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__nand2_1 _06997_ (.A(net64),
    .B(net13),
    .Y(_01217_));
 sky130_fd_sc_hd__nor2_1 _06998_ (.A(_01216_),
    .B(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__xor2_1 _06999_ (.A(_01216_),
    .B(_01217_),
    .X(_01219_));
 sky130_fd_sc_hd__xnor2_1 _07000_ (.A(_01169_),
    .B(_01219_),
    .Y(_01220_));
 sky130_fd_sc_hd__nand2_1 _07001_ (.A(net34),
    .B(net11),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_1 _07002_ (.A(_01220_),
    .B(_01221_),
    .Y(_01222_));
 sky130_fd_sc_hd__xor2_1 _07003_ (.A(_01220_),
    .B(_01221_),
    .X(_01223_));
 sky130_fd_sc_hd__xnor2_1 _07004_ (.A(_01168_),
    .B(_01223_),
    .Y(_01224_));
 sky130_fd_sc_hd__nand2_1 _07005_ (.A(net35),
    .B(net10),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _07006_ (.A(_01224_),
    .B(_01226_),
    .Y(_01227_));
 sky130_fd_sc_hd__xor2_1 _07007_ (.A(_01224_),
    .B(_01226_),
    .X(_01228_));
 sky130_fd_sc_hd__xnor2_1 _07008_ (.A(_01167_),
    .B(_01228_),
    .Y(_01229_));
 sky130_fd_sc_hd__nand2_1 _07009_ (.A(net36),
    .B(net9),
    .Y(_01230_));
 sky130_fd_sc_hd__nor2_1 _07010_ (.A(_01229_),
    .B(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__xor2_1 _07011_ (.A(_01229_),
    .B(_01230_),
    .X(_01232_));
 sky130_fd_sc_hd__xnor2_1 _07012_ (.A(_01166_),
    .B(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__nand2_1 _07013_ (.A(net37),
    .B(net8),
    .Y(_01234_));
 sky130_fd_sc_hd__nor2_1 _07014_ (.A(_01233_),
    .B(_01234_),
    .Y(_01235_));
 sky130_fd_sc_hd__xor2_1 _07015_ (.A(_01233_),
    .B(_01234_),
    .X(_01237_));
 sky130_fd_sc_hd__xnor2_1 _07016_ (.A(_01165_),
    .B(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hd__nand2_1 _07017_ (.A(net38),
    .B(net7),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_1 _07018_ (.A(_01238_),
    .B(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__xor2_1 _07019_ (.A(_01238_),
    .B(_01239_),
    .X(_01241_));
 sky130_fd_sc_hd__xnor2_1 _07020_ (.A(_01164_),
    .B(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__nand2_1 _07021_ (.A(net6),
    .B(net39),
    .Y(_01243_));
 sky130_fd_sc_hd__nor2_1 _07022_ (.A(_01242_),
    .B(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hd__xor2_1 _07023_ (.A(_01242_),
    .B(_01243_),
    .X(_01245_));
 sky130_fd_sc_hd__xnor2_1 _07024_ (.A(_01163_),
    .B(_01245_),
    .Y(_01246_));
 sky130_fd_sc_hd__nand2_1 _07025_ (.A(net5),
    .B(net40),
    .Y(_01248_));
 sky130_fd_sc_hd__nor2_1 _07026_ (.A(_01246_),
    .B(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__xor2_1 _07027_ (.A(_01246_),
    .B(_01248_),
    .X(_01250_));
 sky130_fd_sc_hd__xnor2_1 _07028_ (.A(_01162_),
    .B(_01250_),
    .Y(_01251_));
 sky130_fd_sc_hd__nand2_1 _07029_ (.A(net4),
    .B(net41),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_1 _07030_ (.A(_01251_),
    .B(_01252_),
    .Y(_01253_));
 sky130_fd_sc_hd__xor2_1 _07031_ (.A(_01251_),
    .B(_01252_),
    .X(_01254_));
 sky130_fd_sc_hd__xnor2_1 _07032_ (.A(_01161_),
    .B(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__nand2_1 _07033_ (.A(net3),
    .B(net42),
    .Y(_01256_));
 sky130_fd_sc_hd__nor2_1 _07034_ (.A(_01255_),
    .B(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__xor2_1 _07035_ (.A(_01255_),
    .B(_01256_),
    .X(_01259_));
 sky130_fd_sc_hd__xnor2_1 _07036_ (.A(_01160_),
    .B(_01259_),
    .Y(_01260_));
 sky130_fd_sc_hd__nand2_1 _07037_ (.A(net2),
    .B(net43),
    .Y(_01261_));
 sky130_fd_sc_hd__nor2_1 _07038_ (.A(_01260_),
    .B(_01261_),
    .Y(_01262_));
 sky130_fd_sc_hd__xor2_1 _07039_ (.A(_01260_),
    .B(_01261_),
    .X(_01263_));
 sky130_fd_sc_hd__xnor2_1 _07040_ (.A(_01158_),
    .B(_01263_),
    .Y(_01264_));
 sky130_fd_sc_hd__nand2_1 _07041_ (.A(net32),
    .B(net45),
    .Y(_01265_));
 sky130_fd_sc_hd__nor2_1 _07042_ (.A(_01264_),
    .B(_01265_),
    .Y(_01266_));
 sky130_fd_sc_hd__xor2_1 _07043_ (.A(_01264_),
    .B(_01265_),
    .X(_01267_));
 sky130_fd_sc_hd__xnor2_1 _07044_ (.A(_01157_),
    .B(_01267_),
    .Y(_01268_));
 sky130_fd_sc_hd__nand2_1 _07045_ (.A(net31),
    .B(net46),
    .Y(_01270_));
 sky130_fd_sc_hd__nor2_1 _07046_ (.A(_01268_),
    .B(_01270_),
    .Y(_01271_));
 sky130_fd_sc_hd__xor2_1 _07047_ (.A(_01268_),
    .B(_01270_),
    .X(_01272_));
 sky130_fd_sc_hd__xnor2_1 _07048_ (.A(_01156_),
    .B(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__nand2_1 _07049_ (.A(net30),
    .B(net47),
    .Y(_01274_));
 sky130_fd_sc_hd__nor2_1 _07050_ (.A(_01273_),
    .B(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__xor2_1 _07051_ (.A(_01273_),
    .B(_01274_),
    .X(_01276_));
 sky130_fd_sc_hd__xnor2_1 _07052_ (.A(_01155_),
    .B(_01276_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand2_1 _07053_ (.A(net29),
    .B(net48),
    .Y(_01278_));
 sky130_fd_sc_hd__nor2_1 _07054_ (.A(_01277_),
    .B(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__xor2_1 _07055_ (.A(_01277_),
    .B(_01278_),
    .X(_01281_));
 sky130_fd_sc_hd__xnor2_1 _07056_ (.A(_01154_),
    .B(_01281_),
    .Y(_01282_));
 sky130_fd_sc_hd__nand2_1 _07057_ (.A(net28),
    .B(net49),
    .Y(_01283_));
 sky130_fd_sc_hd__nor2_1 _07058_ (.A(_01282_),
    .B(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__xor2_1 _07059_ (.A(_01282_),
    .B(_01283_),
    .X(_01285_));
 sky130_fd_sc_hd__xnor2_1 _07060_ (.A(_01153_),
    .B(_01285_),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_1 _07061_ (.A(net27),
    .B(net50),
    .Y(_01287_));
 sky130_fd_sc_hd__nor2_1 _07062_ (.A(_01286_),
    .B(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__xor2_1 _07063_ (.A(_01286_),
    .B(_01287_),
    .X(_01289_));
 sky130_fd_sc_hd__xnor2_1 _07064_ (.A(_01152_),
    .B(_01289_),
    .Y(_01290_));
 sky130_fd_sc_hd__nand2_1 _07065_ (.A(net26),
    .B(net51),
    .Y(_01292_));
 sky130_fd_sc_hd__nor2_1 _07066_ (.A(_01290_),
    .B(_01292_),
    .Y(_01293_));
 sky130_fd_sc_hd__xor2_1 _07067_ (.A(_01290_),
    .B(_01292_),
    .X(_01294_));
 sky130_fd_sc_hd__xnor2_1 _07068_ (.A(_01151_),
    .B(_01294_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_1 _07069_ (.A(net23),
    .B(net52),
    .Y(_01296_));
 sky130_fd_sc_hd__nor2_1 _07070_ (.A(_01295_),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__xor2_1 _07071_ (.A(_01295_),
    .B(_01296_),
    .X(_01298_));
 sky130_fd_sc_hd__xnor2_1 _07072_ (.A(_01150_),
    .B(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__nand2_1 _07073_ (.A(net12),
    .B(net53),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_1 _07074_ (.A(_01299_),
    .B(_01300_),
    .Y(_01301_));
 sky130_fd_sc_hd__xor2_1 _07075_ (.A(_01299_),
    .B(_01300_),
    .X(_01303_));
 sky130_fd_sc_hd__xor2_1 _07076_ (.A(_01147_),
    .B(_01303_),
    .X(_01304_));
 sky130_fd_sc_hd__and3_1 _07077_ (.A(net1),
    .B(net54),
    .C(_01304_),
    .X(_01305_));
 sky130_fd_sc_hd__a21oi_1 _07078_ (.A1(net1),
    .A2(net54),
    .B1(_01304_),
    .Y(_01306_));
 sky130_fd_sc_hd__nor2_1 _07079_ (.A(_01305_),
    .B(_01306_),
    .Y(\genblk2[28].rca.ripple_adders[29].fa.sum ));
 sky130_fd_sc_hd__a21o_1 _07080_ (.A1(_01147_),
    .A2(_01303_),
    .B1(_01301_),
    .X(_01307_));
 sky130_fd_sc_hd__a21o_1 _07081_ (.A1(_01150_),
    .A2(_01298_),
    .B1(_01297_),
    .X(_01308_));
 sky130_fd_sc_hd__a21o_1 _07082_ (.A1(_01151_),
    .A2(_01294_),
    .B1(_01293_),
    .X(_01309_));
 sky130_fd_sc_hd__a21o_1 _07083_ (.A1(_01152_),
    .A2(_01289_),
    .B1(_01288_),
    .X(_01310_));
 sky130_fd_sc_hd__a21o_1 _07084_ (.A1(_01153_),
    .A2(_01285_),
    .B1(_01284_),
    .X(_01311_));
 sky130_fd_sc_hd__a21o_1 _07085_ (.A1(_01154_),
    .A2(_01281_),
    .B1(_01279_),
    .X(_01313_));
 sky130_fd_sc_hd__a21o_1 _07086_ (.A1(_01155_),
    .A2(_01276_),
    .B1(_01275_),
    .X(_01314_));
 sky130_fd_sc_hd__a21o_1 _07087_ (.A1(_01156_),
    .A2(_01272_),
    .B1(_01271_),
    .X(_01315_));
 sky130_fd_sc_hd__a21o_1 _07088_ (.A1(_01157_),
    .A2(_01267_),
    .B1(_01266_),
    .X(_01316_));
 sky130_fd_sc_hd__a21o_1 _07089_ (.A1(_01158_),
    .A2(_01263_),
    .B1(_01262_),
    .X(_01317_));
 sky130_fd_sc_hd__a21o_1 _07090_ (.A1(_01160_),
    .A2(_01259_),
    .B1(_01257_),
    .X(_01318_));
 sky130_fd_sc_hd__a21o_1 _07091_ (.A1(_01161_),
    .A2(_01254_),
    .B1(_01253_),
    .X(_01319_));
 sky130_fd_sc_hd__a21o_1 _07092_ (.A1(_01162_),
    .A2(_01250_),
    .B1(_01249_),
    .X(_01320_));
 sky130_fd_sc_hd__a21o_1 _07093_ (.A1(_01163_),
    .A2(_01245_),
    .B1(_01244_),
    .X(_01321_));
 sky130_fd_sc_hd__a21o_1 _07094_ (.A1(_01164_),
    .A2(_01241_),
    .B1(_01240_),
    .X(_01322_));
 sky130_fd_sc_hd__a21o_1 _07095_ (.A1(_01165_),
    .A2(_01237_),
    .B1(_01235_),
    .X(_01324_));
 sky130_fd_sc_hd__a21o_1 _07096_ (.A1(_01166_),
    .A2(_01232_),
    .B1(_01231_),
    .X(_01325_));
 sky130_fd_sc_hd__a21o_1 _07097_ (.A1(_01167_),
    .A2(_01228_),
    .B1(_01227_),
    .X(_01326_));
 sky130_fd_sc_hd__a21o_1 _07098_ (.A1(_01168_),
    .A2(_01223_),
    .B1(_01222_),
    .X(_01327_));
 sky130_fd_sc_hd__a21o_1 _07099_ (.A1(_01169_),
    .A2(_01219_),
    .B1(_01218_),
    .X(_01328_));
 sky130_fd_sc_hd__a21o_1 _07100_ (.A1(_01171_),
    .A2(_01215_),
    .B1(_01213_),
    .X(_01329_));
 sky130_fd_sc_hd__a21o_1 _07101_ (.A1(_01172_),
    .A2(_01210_),
    .B1(_01209_),
    .X(_01330_));
 sky130_fd_sc_hd__a21o_1 _07102_ (.A1(_01173_),
    .A2(_01206_),
    .B1(_01205_),
    .X(_01331_));
 sky130_fd_sc_hd__a21o_1 _07103_ (.A1(_01174_),
    .A2(_01201_),
    .B1(_01200_),
    .X(_01332_));
 sky130_fd_sc_hd__a21o_1 _07104_ (.A1(_01175_),
    .A2(_01197_),
    .B1(_01196_),
    .X(_01333_));
 sky130_fd_sc_hd__a21o_1 _07105_ (.A1(_01176_),
    .A2(_01193_),
    .B1(_01191_),
    .X(_01335_));
 sky130_fd_sc_hd__a21o_1 _07106_ (.A1(_01177_),
    .A2(_01187_),
    .B1(_01186_),
    .X(_01336_));
 sky130_fd_sc_hd__a22o_1 _07107_ (.A1(net44),
    .A2(net22),
    .B1(net24),
    .B2(net33),
    .X(_01337_));
 sky130_fd_sc_hd__nand4_1 _07108_ (.A(net33),
    .B(net44),
    .C(net22),
    .D(net24),
    .Y(_01338_));
 sky130_fd_sc_hd__and2_1 _07109_ (.A(_01337_),
    .B(_01338_),
    .X(_01339_));
 sky130_fd_sc_hd__a21o_1 _07110_ (.A1(_01178_),
    .A2(_01183_),
    .B1(_01179_),
    .X(_01340_));
 sky130_fd_sc_hd__xor2_1 _07111_ (.A(_01339_),
    .B(_01340_),
    .X(_01341_));
 sky130_fd_sc_hd__nand2_1 _07112_ (.A(net55),
    .B(net21),
    .Y(_01342_));
 sky130_fd_sc_hd__and3_1 _07113_ (.A(net55),
    .B(net21),
    .C(_01341_),
    .X(_01343_));
 sky130_fd_sc_hd__nand2b_1 _07114_ (.A_N(_01341_),
    .B(_01342_),
    .Y(_01344_));
 sky130_fd_sc_hd__xor2_1 _07115_ (.A(_01341_),
    .B(_01342_),
    .X(_01346_));
 sky130_fd_sc_hd__xnor2_1 _07116_ (.A(_01336_),
    .B(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__nand2_1 _07117_ (.A(net58),
    .B(net20),
    .Y(_01348_));
 sky130_fd_sc_hd__and3_1 _07118_ (.A(net58),
    .B(net20),
    .C(_01347_),
    .X(_01349_));
 sky130_fd_sc_hd__xnor2_1 _07119_ (.A(_01347_),
    .B(_01348_),
    .Y(_01350_));
 sky130_fd_sc_hd__xor2_1 _07120_ (.A(_01335_),
    .B(_01350_),
    .X(_01351_));
 sky130_fd_sc_hd__nand2_1 _07121_ (.A(net59),
    .B(net19),
    .Y(_01352_));
 sky130_fd_sc_hd__and3_1 _07122_ (.A(net59),
    .B(net19),
    .C(_01351_),
    .X(_01353_));
 sky130_fd_sc_hd__xnor2_1 _07123_ (.A(_01351_),
    .B(_01352_),
    .Y(_01354_));
 sky130_fd_sc_hd__xor2_1 _07124_ (.A(_01333_),
    .B(_01354_),
    .X(_01355_));
 sky130_fd_sc_hd__nand2_1 _07125_ (.A(net60),
    .B(net18),
    .Y(_01357_));
 sky130_fd_sc_hd__and3_1 _07126_ (.A(net60),
    .B(net18),
    .C(_01355_),
    .X(_01358_));
 sky130_fd_sc_hd__xnor2_1 _07127_ (.A(_01355_),
    .B(_01357_),
    .Y(_01359_));
 sky130_fd_sc_hd__xor2_1 _07128_ (.A(_01332_),
    .B(_01359_),
    .X(_01360_));
 sky130_fd_sc_hd__nand2_1 _07129_ (.A(net61),
    .B(net17),
    .Y(_01361_));
 sky130_fd_sc_hd__and3_1 _07130_ (.A(net61),
    .B(net17),
    .C(_01360_),
    .X(_01362_));
 sky130_fd_sc_hd__xnor2_1 _07131_ (.A(_01360_),
    .B(_01361_),
    .Y(_01363_));
 sky130_fd_sc_hd__xnor2_1 _07132_ (.A(_01331_),
    .B(_01363_),
    .Y(_01364_));
 sky130_fd_sc_hd__nand2_1 _07133_ (.A(net62),
    .B(net16),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2_1 _07134_ (.A(_01364_),
    .B(_01365_),
    .Y(_01366_));
 sky130_fd_sc_hd__xor2_1 _07135_ (.A(_01364_),
    .B(_01365_),
    .X(_01368_));
 sky130_fd_sc_hd__xnor2_1 _07136_ (.A(_01330_),
    .B(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hd__nand2_1 _07137_ (.A(net63),
    .B(net15),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_1 _07138_ (.A(_01369_),
    .B(_01370_),
    .Y(_01371_));
 sky130_fd_sc_hd__xor2_1 _07139_ (.A(_01369_),
    .B(_01370_),
    .X(_01372_));
 sky130_fd_sc_hd__xnor2_1 _07140_ (.A(_01329_),
    .B(_01372_),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2_1 _07141_ (.A(net64),
    .B(net14),
    .Y(_01374_));
 sky130_fd_sc_hd__nor2_1 _07142_ (.A(_01373_),
    .B(_01374_),
    .Y(_01375_));
 sky130_fd_sc_hd__xor2_1 _07143_ (.A(_01373_),
    .B(_01374_),
    .X(_01376_));
 sky130_fd_sc_hd__xnor2_1 _07144_ (.A(_01328_),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hd__nand2_1 _07145_ (.A(net34),
    .B(net13),
    .Y(_01379_));
 sky130_fd_sc_hd__nor2_1 _07146_ (.A(_01377_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__xor2_1 _07147_ (.A(_01377_),
    .B(_01379_),
    .X(_01381_));
 sky130_fd_sc_hd__xnor2_1 _07148_ (.A(_01327_),
    .B(_01381_),
    .Y(_01382_));
 sky130_fd_sc_hd__nand2_1 _07149_ (.A(net35),
    .B(net11),
    .Y(_01383_));
 sky130_fd_sc_hd__nor2_1 _07150_ (.A(_01382_),
    .B(_01383_),
    .Y(_01384_));
 sky130_fd_sc_hd__xor2_1 _07151_ (.A(_01382_),
    .B(_01383_),
    .X(_01385_));
 sky130_fd_sc_hd__xnor2_1 _07152_ (.A(_01326_),
    .B(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hd__nand2_1 _07153_ (.A(net36),
    .B(net10),
    .Y(_01387_));
 sky130_fd_sc_hd__nor2_1 _07154_ (.A(_01386_),
    .B(_01387_),
    .Y(_01388_));
 sky130_fd_sc_hd__xor2_1 _07155_ (.A(_01386_),
    .B(_01387_),
    .X(_01390_));
 sky130_fd_sc_hd__xnor2_1 _07156_ (.A(_01325_),
    .B(_01390_),
    .Y(_01391_));
 sky130_fd_sc_hd__nand2_1 _07157_ (.A(net37),
    .B(net9),
    .Y(_01392_));
 sky130_fd_sc_hd__nor2_1 _07158_ (.A(_01391_),
    .B(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__xor2_1 _07159_ (.A(_01391_),
    .B(_01392_),
    .X(_01394_));
 sky130_fd_sc_hd__xnor2_1 _07160_ (.A(_01324_),
    .B(_01394_),
    .Y(_01395_));
 sky130_fd_sc_hd__nand2_1 _07161_ (.A(net38),
    .B(net8),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_1 _07162_ (.A(_01395_),
    .B(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hd__xor2_1 _07163_ (.A(_01395_),
    .B(_01396_),
    .X(_01398_));
 sky130_fd_sc_hd__xnor2_1 _07164_ (.A(_01322_),
    .B(_01398_),
    .Y(_01399_));
 sky130_fd_sc_hd__nand2_1 _07165_ (.A(net7),
    .B(net39),
    .Y(_01401_));
 sky130_fd_sc_hd__nor2_1 _07166_ (.A(_01399_),
    .B(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__xor2_1 _07167_ (.A(_01399_),
    .B(_01401_),
    .X(_01403_));
 sky130_fd_sc_hd__xnor2_1 _07168_ (.A(_01321_),
    .B(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__nand2_1 _07169_ (.A(net6),
    .B(net40),
    .Y(_01405_));
 sky130_fd_sc_hd__nor2_1 _07170_ (.A(_01404_),
    .B(_01405_),
    .Y(_01406_));
 sky130_fd_sc_hd__xor2_1 _07171_ (.A(_01404_),
    .B(_01405_),
    .X(_01407_));
 sky130_fd_sc_hd__xnor2_1 _07172_ (.A(_01320_),
    .B(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__nand2_1 _07173_ (.A(net5),
    .B(net41),
    .Y(_01409_));
 sky130_fd_sc_hd__nor2_1 _07174_ (.A(_01408_),
    .B(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__xor2_1 _07175_ (.A(_01408_),
    .B(_01409_),
    .X(_01412_));
 sky130_fd_sc_hd__xnor2_1 _07176_ (.A(_01319_),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__nand2_1 _07177_ (.A(net4),
    .B(net42),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_1 _07178_ (.A(_01413_),
    .B(_01414_),
    .Y(_01415_));
 sky130_fd_sc_hd__xor2_1 _07179_ (.A(_01413_),
    .B(_01414_),
    .X(_01416_));
 sky130_fd_sc_hd__xnor2_1 _07180_ (.A(_01318_),
    .B(_01416_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2_1 _07181_ (.A(net3),
    .B(net43),
    .Y(_01418_));
 sky130_fd_sc_hd__nor2_1 _07182_ (.A(_01417_),
    .B(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__xor2_1 _07183_ (.A(_01417_),
    .B(_01418_),
    .X(_01420_));
 sky130_fd_sc_hd__xnor2_1 _07184_ (.A(_01317_),
    .B(_01420_),
    .Y(_01421_));
 sky130_fd_sc_hd__nand2_1 _07185_ (.A(net2),
    .B(net45),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_1 _07186_ (.A(_01421_),
    .B(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__xor2_1 _07187_ (.A(_01421_),
    .B(_01423_),
    .X(_01425_));
 sky130_fd_sc_hd__xnor2_1 _07188_ (.A(_01316_),
    .B(_01425_),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_1 _07189_ (.A(net32),
    .B(net46),
    .Y(_01427_));
 sky130_fd_sc_hd__nor2_1 _07190_ (.A(_01426_),
    .B(_01427_),
    .Y(_01428_));
 sky130_fd_sc_hd__xor2_1 _07191_ (.A(_01426_),
    .B(_01427_),
    .X(_01429_));
 sky130_fd_sc_hd__xnor2_1 _07192_ (.A(_01315_),
    .B(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__nand2_1 _07193_ (.A(net31),
    .B(net47),
    .Y(_01431_));
 sky130_fd_sc_hd__nor2_1 _07194_ (.A(_01430_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__xor2_1 _07195_ (.A(_01430_),
    .B(_01431_),
    .X(_01434_));
 sky130_fd_sc_hd__xnor2_1 _07196_ (.A(_01314_),
    .B(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2_1 _07197_ (.A(net30),
    .B(net48),
    .Y(_01436_));
 sky130_fd_sc_hd__nor2_1 _07198_ (.A(_01435_),
    .B(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__xor2_1 _07199_ (.A(_01435_),
    .B(_01436_),
    .X(_01438_));
 sky130_fd_sc_hd__xnor2_1 _07200_ (.A(_01313_),
    .B(_01438_),
    .Y(_01439_));
 sky130_fd_sc_hd__nand2_1 _07201_ (.A(net29),
    .B(net49),
    .Y(_01440_));
 sky130_fd_sc_hd__nor2_1 _07202_ (.A(_01439_),
    .B(_01440_),
    .Y(_01441_));
 sky130_fd_sc_hd__xor2_1 _07203_ (.A(_01439_),
    .B(_01440_),
    .X(_01442_));
 sky130_fd_sc_hd__xnor2_1 _07204_ (.A(_01311_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__nand2_1 _07205_ (.A(net28),
    .B(net50),
    .Y(_01445_));
 sky130_fd_sc_hd__nor2_1 _07206_ (.A(_01443_),
    .B(_01445_),
    .Y(_01446_));
 sky130_fd_sc_hd__xor2_1 _07207_ (.A(_01443_),
    .B(_01445_),
    .X(_01447_));
 sky130_fd_sc_hd__xnor2_1 _07208_ (.A(_01310_),
    .B(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__nand2_1 _07209_ (.A(net27),
    .B(net51),
    .Y(_01449_));
 sky130_fd_sc_hd__nor2_1 _07210_ (.A(_01448_),
    .B(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__xor2_1 _07211_ (.A(_01448_),
    .B(_01449_),
    .X(_01451_));
 sky130_fd_sc_hd__xnor2_1 _07212_ (.A(_01309_),
    .B(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__nand2_1 _07213_ (.A(net26),
    .B(net52),
    .Y(_01453_));
 sky130_fd_sc_hd__nor2_1 _07214_ (.A(_01452_),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__xor2_1 _07215_ (.A(_01452_),
    .B(_01453_),
    .X(_01456_));
 sky130_fd_sc_hd__xnor2_1 _07216_ (.A(_01308_),
    .B(_01456_),
    .Y(_01457_));
 sky130_fd_sc_hd__nand2_1 _07217_ (.A(net23),
    .B(net53),
    .Y(_01458_));
 sky130_fd_sc_hd__nor2_1 _07218_ (.A(_01457_),
    .B(_01458_),
    .Y(_01459_));
 sky130_fd_sc_hd__xor2_1 _07219_ (.A(_01457_),
    .B(_01458_),
    .X(_01460_));
 sky130_fd_sc_hd__xnor2_1 _07220_ (.A(_01307_),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__nand2_1 _07221_ (.A(net12),
    .B(net54),
    .Y(_01462_));
 sky130_fd_sc_hd__nor2_1 _07222_ (.A(_01461_),
    .B(_01462_),
    .Y(_01463_));
 sky130_fd_sc_hd__xor2_1 _07223_ (.A(_01461_),
    .B(_01462_),
    .X(_01464_));
 sky130_fd_sc_hd__xor2_1 _07224_ (.A(_01305_),
    .B(_01464_),
    .X(_01465_));
 sky130_fd_sc_hd__and3_1 _07225_ (.A(net1),
    .B(net56),
    .C(_01465_),
    .X(_01467_));
 sky130_fd_sc_hd__a21oi_1 _07226_ (.A1(net1),
    .A2(net56),
    .B1(_01465_),
    .Y(_01468_));
 sky130_fd_sc_hd__nor2_1 _07227_ (.A(_01467_),
    .B(_01468_),
    .Y(\genblk2[29].rca.ripple_adders[30].fa.sum ));
 sky130_fd_sc_hd__nand2_1 _07228_ (.A(net12),
    .B(net56),
    .Y(_01469_));
 sky130_fd_sc_hd__a21o_1 _07229_ (.A1(_01305_),
    .A2(_01464_),
    .B1(_01463_),
    .X(_01470_));
 sky130_fd_sc_hd__nand2_1 _07230_ (.A(net23),
    .B(net54),
    .Y(_01471_));
 sky130_fd_sc_hd__a21o_1 _07231_ (.A1(_01307_),
    .A2(_01460_),
    .B1(_01459_),
    .X(_01472_));
 sky130_fd_sc_hd__nand2_1 _07232_ (.A(net26),
    .B(net53),
    .Y(_01473_));
 sky130_fd_sc_hd__a21o_1 _07233_ (.A1(_01308_),
    .A2(_01456_),
    .B1(_01454_),
    .X(_01474_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(net27),
    .B(net52),
    .Y(_01475_));
 sky130_fd_sc_hd__a21o_1 _07235_ (.A1(_01309_),
    .A2(_01451_),
    .B1(_01450_),
    .X(_01477_));
 sky130_fd_sc_hd__nand2_1 _07236_ (.A(net28),
    .B(net51),
    .Y(_01478_));
 sky130_fd_sc_hd__a21o_1 _07237_ (.A1(_01310_),
    .A2(_01447_),
    .B1(_01446_),
    .X(_01479_));
 sky130_fd_sc_hd__nand2_1 _07238_ (.A(net29),
    .B(net50),
    .Y(_01480_));
 sky130_fd_sc_hd__a21o_1 _07239_ (.A1(_01311_),
    .A2(_01442_),
    .B1(_01441_),
    .X(_01481_));
 sky130_fd_sc_hd__nand2_1 _07240_ (.A(net30),
    .B(net49),
    .Y(_01482_));
 sky130_fd_sc_hd__a21o_1 _07241_ (.A1(_01313_),
    .A2(_01438_),
    .B1(_01437_),
    .X(_01483_));
 sky130_fd_sc_hd__nand2_1 _07242_ (.A(net31),
    .B(net48),
    .Y(_01484_));
 sky130_fd_sc_hd__a21o_1 _07243_ (.A1(_01314_),
    .A2(_01434_),
    .B1(_01432_),
    .X(_01485_));
 sky130_fd_sc_hd__nand2_1 _07244_ (.A(net32),
    .B(net47),
    .Y(_01486_));
 sky130_fd_sc_hd__a21o_1 _07245_ (.A1(_01315_),
    .A2(_01429_),
    .B1(_01428_),
    .X(_01488_));
 sky130_fd_sc_hd__nand2_1 _07246_ (.A(net2),
    .B(net46),
    .Y(_01489_));
 sky130_fd_sc_hd__a21o_1 _07247_ (.A1(_01316_),
    .A2(_01425_),
    .B1(_01424_),
    .X(_01490_));
 sky130_fd_sc_hd__nand2_1 _07248_ (.A(net3),
    .B(net45),
    .Y(_01491_));
 sky130_fd_sc_hd__a21o_1 _07249_ (.A1(_01317_),
    .A2(_01420_),
    .B1(_01419_),
    .X(_01492_));
 sky130_fd_sc_hd__nand2_1 _07250_ (.A(net4),
    .B(net43),
    .Y(_01493_));
 sky130_fd_sc_hd__a21o_1 _07251_ (.A1(_01318_),
    .A2(_01416_),
    .B1(_01415_),
    .X(_01494_));
 sky130_fd_sc_hd__nand2_1 _07252_ (.A(net5),
    .B(net42),
    .Y(_01495_));
 sky130_fd_sc_hd__a21o_1 _07253_ (.A1(_01319_),
    .A2(_01412_),
    .B1(_01410_),
    .X(_01496_));
 sky130_fd_sc_hd__nand2_1 _07254_ (.A(net6),
    .B(net41),
    .Y(_01497_));
 sky130_fd_sc_hd__a21o_1 _07255_ (.A1(_01320_),
    .A2(_01407_),
    .B1(_01406_),
    .X(_01499_));
 sky130_fd_sc_hd__nand2_1 _07256_ (.A(net7),
    .B(net40),
    .Y(_01500_));
 sky130_fd_sc_hd__a21o_1 _07257_ (.A1(_01321_),
    .A2(_01403_),
    .B1(_01402_),
    .X(_01501_));
 sky130_fd_sc_hd__nand2_1 _07258_ (.A(net39),
    .B(net8),
    .Y(_01502_));
 sky130_fd_sc_hd__a21o_1 _07259_ (.A1(_01322_),
    .A2(_01398_),
    .B1(_01397_),
    .X(_01503_));
 sky130_fd_sc_hd__nand2_1 _07260_ (.A(net38),
    .B(net9),
    .Y(_01504_));
 sky130_fd_sc_hd__a21o_1 _07261_ (.A1(_01324_),
    .A2(_01394_),
    .B1(_01393_),
    .X(_01505_));
 sky130_fd_sc_hd__nand2_1 _07262_ (.A(net37),
    .B(net10),
    .Y(_01506_));
 sky130_fd_sc_hd__a21o_1 _07263_ (.A1(_01325_),
    .A2(_01390_),
    .B1(_01388_),
    .X(_01507_));
 sky130_fd_sc_hd__nand2_1 _07264_ (.A(net36),
    .B(net11),
    .Y(_01508_));
 sky130_fd_sc_hd__a21o_1 _07265_ (.A1(_01326_),
    .A2(_01385_),
    .B1(_01384_),
    .X(_01510_));
 sky130_fd_sc_hd__nand2_1 _07266_ (.A(net35),
    .B(net13),
    .Y(_01511_));
 sky130_fd_sc_hd__a21o_1 _07267_ (.A1(_01327_),
    .A2(_01381_),
    .B1(_01380_),
    .X(_01512_));
 sky130_fd_sc_hd__nand2_1 _07268_ (.A(net34),
    .B(net14),
    .Y(_01513_));
 sky130_fd_sc_hd__a21o_1 _07269_ (.A1(_01328_),
    .A2(_01376_),
    .B1(_01375_),
    .X(_01514_));
 sky130_fd_sc_hd__nand2_1 _07270_ (.A(net64),
    .B(net15),
    .Y(_01515_));
 sky130_fd_sc_hd__a21o_1 _07271_ (.A1(_01329_),
    .A2(_01372_),
    .B1(_01371_),
    .X(_01516_));
 sky130_fd_sc_hd__nand2_1 _07272_ (.A(net63),
    .B(net16),
    .Y(_01517_));
 sky130_fd_sc_hd__a21o_1 _07273_ (.A1(_01330_),
    .A2(_01368_),
    .B1(_01366_),
    .X(_01518_));
 sky130_fd_sc_hd__nand2_1 _07274_ (.A(net62),
    .B(net17),
    .Y(_01519_));
 sky130_fd_sc_hd__a21o_1 _07275_ (.A1(_01331_),
    .A2(_01363_),
    .B1(_01362_),
    .X(_01521_));
 sky130_fd_sc_hd__nand2_1 _07276_ (.A(net61),
    .B(net18),
    .Y(_01522_));
 sky130_fd_sc_hd__a21o_1 _07277_ (.A1(_01332_),
    .A2(_01359_),
    .B1(_01358_),
    .X(_01523_));
 sky130_fd_sc_hd__nand2_1 _07278_ (.A(net60),
    .B(net19),
    .Y(_01524_));
 sky130_fd_sc_hd__a21o_1 _07279_ (.A1(_01333_),
    .A2(_01354_),
    .B1(_01353_),
    .X(_01525_));
 sky130_fd_sc_hd__nand2_1 _07280_ (.A(net59),
    .B(net20),
    .Y(_01526_));
 sky130_fd_sc_hd__a21o_1 _07281_ (.A1(_01335_),
    .A2(_01350_),
    .B1(_01349_),
    .X(_01527_));
 sky130_fd_sc_hd__nand2_1 _07282_ (.A(net58),
    .B(net21),
    .Y(_01528_));
 sky130_fd_sc_hd__a21o_1 _07283_ (.A1(_01336_),
    .A2(_01344_),
    .B1(_01343_),
    .X(_01529_));
 sky130_fd_sc_hd__nand2_1 _07284_ (.A(net55),
    .B(net22),
    .Y(_01530_));
 sky130_fd_sc_hd__a21boi_1 _07285_ (.A1(_01337_),
    .A2(_01340_),
    .B1_N(_01338_),
    .Y(_01532_));
 sky130_fd_sc_hd__a22o_1 _07286_ (.A1(net44),
    .A2(net24),
    .B1(net25),
    .B2(net33),
    .X(_01533_));
 sky130_fd_sc_hd__and3_1 _07287_ (.A(net33),
    .B(net24),
    .C(net25),
    .X(_01534_));
 sky130_fd_sc_hd__a21bo_1 _07288_ (.A1(net44),
    .A2(_01534_),
    .B1_N(_01533_),
    .X(_01535_));
 sky130_fd_sc_hd__nor2_1 _07289_ (.A(_01532_),
    .B(_01535_),
    .Y(_01536_));
 sky130_fd_sc_hd__xor2_1 _07290_ (.A(_01532_),
    .B(_01535_),
    .X(_01537_));
 sky130_fd_sc_hd__and3_1 _07291_ (.A(net55),
    .B(net22),
    .C(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__xnor2_1 _07292_ (.A(_01530_),
    .B(_01537_),
    .Y(_01539_));
 sky130_fd_sc_hd__xor2_1 _07293_ (.A(_01529_),
    .B(_01539_),
    .X(_01540_));
 sky130_fd_sc_hd__and3_1 _07294_ (.A(net58),
    .B(net21),
    .C(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__xnor2_1 _07295_ (.A(_01528_),
    .B(_01540_),
    .Y(_01543_));
 sky130_fd_sc_hd__xor2_1 _07296_ (.A(_01527_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__and3_1 _07297_ (.A(net59),
    .B(net20),
    .C(_01544_),
    .X(_01545_));
 sky130_fd_sc_hd__xnor2_1 _07298_ (.A(_01526_),
    .B(_01544_),
    .Y(_01546_));
 sky130_fd_sc_hd__xor2_1 _07299_ (.A(_01525_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__and3_1 _07300_ (.A(net60),
    .B(net19),
    .C(_01547_),
    .X(_01548_));
 sky130_fd_sc_hd__xnor2_1 _07301_ (.A(_01524_),
    .B(_01547_),
    .Y(_01549_));
 sky130_fd_sc_hd__xor2_1 _07302_ (.A(_01523_),
    .B(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__and3_1 _07303_ (.A(net61),
    .B(net18),
    .C(_01550_),
    .X(_01551_));
 sky130_fd_sc_hd__xnor2_1 _07304_ (.A(_01522_),
    .B(_01550_),
    .Y(_01552_));
 sky130_fd_sc_hd__xor2_1 _07305_ (.A(_01521_),
    .B(_01552_),
    .X(_01554_));
 sky130_fd_sc_hd__and3_1 _07306_ (.A(net62),
    .B(net17),
    .C(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__xnor2_1 _07307_ (.A(_01519_),
    .B(_01554_),
    .Y(_01556_));
 sky130_fd_sc_hd__xor2_1 _07308_ (.A(_01518_),
    .B(_01556_),
    .X(_01557_));
 sky130_fd_sc_hd__and3_1 _07309_ (.A(net63),
    .B(net16),
    .C(_01557_),
    .X(_01558_));
 sky130_fd_sc_hd__xnor2_1 _07310_ (.A(_01517_),
    .B(_01557_),
    .Y(_01559_));
 sky130_fd_sc_hd__xor2_1 _07311_ (.A(_01516_),
    .B(_01559_),
    .X(_01560_));
 sky130_fd_sc_hd__and3_1 _07312_ (.A(net64),
    .B(net15),
    .C(_01560_),
    .X(_01561_));
 sky130_fd_sc_hd__xnor2_1 _07313_ (.A(_01515_),
    .B(_01560_),
    .Y(_01562_));
 sky130_fd_sc_hd__xor2_1 _07314_ (.A(_01514_),
    .B(_01562_),
    .X(_01563_));
 sky130_fd_sc_hd__and3_1 _07315_ (.A(net34),
    .B(net14),
    .C(_01563_),
    .X(_01565_));
 sky130_fd_sc_hd__xnor2_1 _07316_ (.A(_01513_),
    .B(_01563_),
    .Y(_01566_));
 sky130_fd_sc_hd__xor2_1 _07317_ (.A(_01512_),
    .B(_01566_),
    .X(_01567_));
 sky130_fd_sc_hd__and3_1 _07318_ (.A(net35),
    .B(net13),
    .C(_01567_),
    .X(_01568_));
 sky130_fd_sc_hd__xnor2_1 _07319_ (.A(_01511_),
    .B(_01567_),
    .Y(_01569_));
 sky130_fd_sc_hd__xor2_1 _07320_ (.A(_01510_),
    .B(_01569_),
    .X(_01570_));
 sky130_fd_sc_hd__and3_1 _07321_ (.A(net36),
    .B(net11),
    .C(_01570_),
    .X(_01571_));
 sky130_fd_sc_hd__xnor2_1 _07322_ (.A(_01508_),
    .B(_01570_),
    .Y(_01572_));
 sky130_fd_sc_hd__xor2_1 _07323_ (.A(_01507_),
    .B(_01572_),
    .X(_01573_));
 sky130_fd_sc_hd__and3_1 _07324_ (.A(net37),
    .B(net10),
    .C(_01573_),
    .X(_01574_));
 sky130_fd_sc_hd__xnor2_1 _07325_ (.A(_01506_),
    .B(_01573_),
    .Y(_01576_));
 sky130_fd_sc_hd__xor2_1 _07326_ (.A(_01505_),
    .B(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__and3_1 _07327_ (.A(net38),
    .B(net9),
    .C(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__xnor2_1 _07328_ (.A(_01504_),
    .B(_01577_),
    .Y(_01579_));
 sky130_fd_sc_hd__xor2_1 _07329_ (.A(_01503_),
    .B(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__and3_1 _07330_ (.A(net39),
    .B(net8),
    .C(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__xnor2_1 _07331_ (.A(_01502_),
    .B(_01580_),
    .Y(_01582_));
 sky130_fd_sc_hd__xor2_1 _07332_ (.A(_01501_),
    .B(_01582_),
    .X(_01583_));
 sky130_fd_sc_hd__and3_1 _07333_ (.A(net7),
    .B(net40),
    .C(_01583_),
    .X(_01584_));
 sky130_fd_sc_hd__xnor2_1 _07334_ (.A(_01500_),
    .B(_01583_),
    .Y(_01585_));
 sky130_fd_sc_hd__xor2_1 _07335_ (.A(_01499_),
    .B(_01585_),
    .X(_01587_));
 sky130_fd_sc_hd__and3_1 _07336_ (.A(net6),
    .B(net41),
    .C(_01587_),
    .X(_01588_));
 sky130_fd_sc_hd__xnor2_1 _07337_ (.A(_01497_),
    .B(_01587_),
    .Y(_01589_));
 sky130_fd_sc_hd__xor2_1 _07338_ (.A(_01496_),
    .B(_01589_),
    .X(_01590_));
 sky130_fd_sc_hd__and3_1 _07339_ (.A(net5),
    .B(net42),
    .C(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__xnor2_1 _07340_ (.A(_01495_),
    .B(_01590_),
    .Y(_01592_));
 sky130_fd_sc_hd__xor2_1 _07341_ (.A(_01494_),
    .B(_01592_),
    .X(_01593_));
 sky130_fd_sc_hd__and3_1 _07342_ (.A(net4),
    .B(net43),
    .C(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__xnor2_1 _07343_ (.A(_01493_),
    .B(_01593_),
    .Y(_01595_));
 sky130_fd_sc_hd__xor2_1 _07344_ (.A(_01492_),
    .B(_01595_),
    .X(_01596_));
 sky130_fd_sc_hd__and3_1 _07345_ (.A(net3),
    .B(net45),
    .C(_01596_),
    .X(_01598_));
 sky130_fd_sc_hd__xnor2_1 _07346_ (.A(_01491_),
    .B(_01596_),
    .Y(_01599_));
 sky130_fd_sc_hd__xor2_1 _07347_ (.A(_01490_),
    .B(_01599_),
    .X(_01600_));
 sky130_fd_sc_hd__and3_1 _07348_ (.A(net2),
    .B(net46),
    .C(_01600_),
    .X(_01601_));
 sky130_fd_sc_hd__xnor2_1 _07349_ (.A(_01489_),
    .B(_01600_),
    .Y(_01602_));
 sky130_fd_sc_hd__xor2_1 _07350_ (.A(_01488_),
    .B(_01602_),
    .X(_01603_));
 sky130_fd_sc_hd__and3_1 _07351_ (.A(net32),
    .B(net47),
    .C(_01603_),
    .X(_01604_));
 sky130_fd_sc_hd__xnor2_1 _07352_ (.A(_01486_),
    .B(_01603_),
    .Y(_01605_));
 sky130_fd_sc_hd__xor2_1 _07353_ (.A(_01485_),
    .B(_01605_),
    .X(_01606_));
 sky130_fd_sc_hd__and3_1 _07354_ (.A(net31),
    .B(net48),
    .C(_01606_),
    .X(_01607_));
 sky130_fd_sc_hd__xnor2_1 _07355_ (.A(_01484_),
    .B(_01606_),
    .Y(_01609_));
 sky130_fd_sc_hd__xor2_1 _07356_ (.A(_01483_),
    .B(_01609_),
    .X(_01610_));
 sky130_fd_sc_hd__and3_1 _07357_ (.A(net30),
    .B(net49),
    .C(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__xnor2_1 _07358_ (.A(_01482_),
    .B(_01610_),
    .Y(_01612_));
 sky130_fd_sc_hd__xor2_1 _07359_ (.A(_01481_),
    .B(_01612_),
    .X(_01613_));
 sky130_fd_sc_hd__and3_1 _07360_ (.A(net29),
    .B(net50),
    .C(_01613_),
    .X(_01614_));
 sky130_fd_sc_hd__xnor2_1 _07361_ (.A(_01480_),
    .B(_01613_),
    .Y(_01615_));
 sky130_fd_sc_hd__xor2_1 _07362_ (.A(_01479_),
    .B(_01615_),
    .X(_01616_));
 sky130_fd_sc_hd__and3_1 _07363_ (.A(net28),
    .B(net51),
    .C(_01616_),
    .X(_01617_));
 sky130_fd_sc_hd__xnor2_1 _07364_ (.A(_01478_),
    .B(_01616_),
    .Y(_01618_));
 sky130_fd_sc_hd__xor2_1 _07365_ (.A(_01477_),
    .B(_01618_),
    .X(_01620_));
 sky130_fd_sc_hd__and3_1 _07366_ (.A(net27),
    .B(net52),
    .C(_01620_),
    .X(_01621_));
 sky130_fd_sc_hd__xnor2_1 _07367_ (.A(_01475_),
    .B(_01620_),
    .Y(_01622_));
 sky130_fd_sc_hd__xor2_1 _07368_ (.A(_01474_),
    .B(_01622_),
    .X(_01623_));
 sky130_fd_sc_hd__and3_1 _07369_ (.A(net26),
    .B(net53),
    .C(_01623_),
    .X(_01624_));
 sky130_fd_sc_hd__xnor2_1 _07370_ (.A(_01473_),
    .B(_01623_),
    .Y(_01625_));
 sky130_fd_sc_hd__xor2_1 _07371_ (.A(_01472_),
    .B(_01625_),
    .X(_01626_));
 sky130_fd_sc_hd__and3_1 _07372_ (.A(net23),
    .B(net54),
    .C(_01626_),
    .X(_01627_));
 sky130_fd_sc_hd__xnor2_1 _07373_ (.A(_01471_),
    .B(_01626_),
    .Y(_01628_));
 sky130_fd_sc_hd__xor2_1 _07374_ (.A(_01470_),
    .B(_01628_),
    .X(_01629_));
 sky130_fd_sc_hd__and3_1 _07375_ (.A(net12),
    .B(net56),
    .C(_01629_),
    .X(_01631_));
 sky130_fd_sc_hd__xnor2_1 _07376_ (.A(_01469_),
    .B(_01629_),
    .Y(_01632_));
 sky130_fd_sc_hd__xor2_1 _07377_ (.A(_01467_),
    .B(_01632_),
    .X(_01633_));
 sky130_fd_sc_hd__and3_1 _07378_ (.A(net1),
    .B(net57),
    .C(_01633_),
    .X(_01634_));
 sky130_fd_sc_hd__a21oi_1 _07379_ (.A1(net1),
    .A2(net57),
    .B1(_01633_),
    .Y(_01635_));
 sky130_fd_sc_hd__nor2_1 _07380_ (.A(_01634_),
    .B(_01635_),
    .Y(\genblk2[30].rca.ripple_adders[31].fa.sum ));
 sky130_fd_sc_hd__a21oi_1 _07381_ (.A1(_01529_),
    .A2(_01539_),
    .B1(_01538_),
    .Y(_01636_));
 sky130_fd_sc_hd__or2_1 _07382_ (.A(net33),
    .B(net44),
    .X(_01637_));
 sky130_fd_sc_hd__o211a_1 _07383_ (.A1(net24),
    .A2(_00384_),
    .B1(_01637_),
    .C1(net25),
    .X(_01638_));
 sky130_fd_sc_hd__o211a_1 _07384_ (.A1(_01536_),
    .A2(_01638_),
    .B1(net55),
    .C1(net24),
    .X(_01639_));
 sky130_fd_sc_hd__a211oi_1 _07385_ (.A1(net55),
    .A2(net24),
    .B1(_01536_),
    .C1(_01638_),
    .Y(_01641_));
 sky130_fd_sc_hd__nor2_1 _07386_ (.A(_01639_),
    .B(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__and2b_1 _07387_ (.A_N(_01636_),
    .B(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__xnor2_1 _07388_ (.A(_01636_),
    .B(_01642_),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _07389_ (.A(net58),
    .B(net22),
    .Y(_01645_));
 sky130_fd_sc_hd__and3_1 _07390_ (.A(net58),
    .B(net22),
    .C(_01644_),
    .X(_01646_));
 sky130_fd_sc_hd__a21o_1 _07391_ (.A1(_01527_),
    .A2(_01543_),
    .B1(_01541_),
    .X(_01647_));
 sky130_fd_sc_hd__xnor2_1 _07392_ (.A(_01644_),
    .B(_01645_),
    .Y(_01648_));
 sky130_fd_sc_hd__a21oi_1 _07393_ (.A1(_01647_),
    .A2(_01648_),
    .B1(_01646_),
    .Y(_01649_));
 sky130_fd_sc_hd__or2_1 _07394_ (.A(net55),
    .B(_01637_),
    .X(_01650_));
 sky130_fd_sc_hd__nand2_1 _07395_ (.A(net55),
    .B(_01637_),
    .Y(_01652_));
 sky130_fd_sc_hd__a311o_1 _07396_ (.A1(net25),
    .A2(_01650_),
    .A3(_01652_),
    .B1(_01639_),
    .C1(_01643_),
    .X(_01653_));
 sky130_fd_sc_hd__nand2_1 _07397_ (.A(net58),
    .B(net24),
    .Y(_01654_));
 sky130_fd_sc_hd__nand2b_1 _07398_ (.A_N(_01654_),
    .B(_01653_),
    .Y(_01655_));
 sky130_fd_sc_hd__xnor2_1 _07399_ (.A(_01653_),
    .B(_01654_),
    .Y(_01656_));
 sky130_fd_sc_hd__nand2b_1 _07400_ (.A_N(_01649_),
    .B(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__xnor2_1 _07401_ (.A(_01649_),
    .B(_01656_),
    .Y(_01658_));
 sky130_fd_sc_hd__nand2_1 _07402_ (.A(net59),
    .B(net22),
    .Y(_01659_));
 sky130_fd_sc_hd__and3_1 _07403_ (.A(net59),
    .B(net22),
    .C(_01658_),
    .X(_01660_));
 sky130_fd_sc_hd__xor2_1 _07404_ (.A(_01647_),
    .B(_01648_),
    .X(_01661_));
 sky130_fd_sc_hd__nand2_1 _07405_ (.A(net59),
    .B(net21),
    .Y(_01663_));
 sky130_fd_sc_hd__and3_1 _07406_ (.A(net59),
    .B(net21),
    .C(_01661_),
    .X(_01664_));
 sky130_fd_sc_hd__a21o_1 _07407_ (.A1(_01525_),
    .A2(_01546_),
    .B1(_01545_),
    .X(_01665_));
 sky130_fd_sc_hd__xnor2_1 _07408_ (.A(_01661_),
    .B(_01663_),
    .Y(_01666_));
 sky130_fd_sc_hd__a21o_1 _07409_ (.A1(_01665_),
    .A2(_01666_),
    .B1(_01664_),
    .X(_01667_));
 sky130_fd_sc_hd__xnor2_1 _07410_ (.A(_01658_),
    .B(_01659_),
    .Y(_01668_));
 sky130_fd_sc_hd__a21oi_1 _07411_ (.A1(_01667_),
    .A2(_01668_),
    .B1(_01660_),
    .Y(_01669_));
 sky130_fd_sc_hd__nand2_1 _07412_ (.A(net59),
    .B(net24),
    .Y(_01670_));
 sky130_fd_sc_hd__o21a_1 _07413_ (.A1(net58),
    .A2(_01650_),
    .B1(net25),
    .X(_01671_));
 sky130_fd_sc_hd__a21bo_1 _07414_ (.A1(net58),
    .A2(_01650_),
    .B1_N(_01671_),
    .X(_01672_));
 sky130_fd_sc_hd__and3_1 _07415_ (.A(_01655_),
    .B(_01657_),
    .C(_01672_),
    .X(_01674_));
 sky130_fd_sc_hd__nor2_1 _07416_ (.A(_01670_),
    .B(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__xnor2_1 _07417_ (.A(_01670_),
    .B(_01674_),
    .Y(_01676_));
 sky130_fd_sc_hd__nor2_1 _07418_ (.A(_01669_),
    .B(_01676_),
    .Y(_01677_));
 sky130_fd_sc_hd__xor2_1 _07419_ (.A(_01669_),
    .B(_01676_),
    .X(_01678_));
 sky130_fd_sc_hd__nand2_1 _07420_ (.A(net60),
    .B(net22),
    .Y(_01679_));
 sky130_fd_sc_hd__and3_1 _07421_ (.A(net60),
    .B(net22),
    .C(_01678_),
    .X(_01680_));
 sky130_fd_sc_hd__xor2_1 _07422_ (.A(_01667_),
    .B(_01668_),
    .X(_01681_));
 sky130_fd_sc_hd__nand2_1 _07423_ (.A(net60),
    .B(net21),
    .Y(_01682_));
 sky130_fd_sc_hd__and3_1 _07424_ (.A(net60),
    .B(net21),
    .C(_01681_),
    .X(_01683_));
 sky130_fd_sc_hd__xor2_1 _07425_ (.A(_01665_),
    .B(_01666_),
    .X(_01685_));
 sky130_fd_sc_hd__nand2_1 _07426_ (.A(net60),
    .B(net20),
    .Y(_01686_));
 sky130_fd_sc_hd__and3_1 _07427_ (.A(net60),
    .B(net20),
    .C(_01685_),
    .X(_01687_));
 sky130_fd_sc_hd__a21o_1 _07428_ (.A1(_01523_),
    .A2(_01549_),
    .B1(_01548_),
    .X(_01688_));
 sky130_fd_sc_hd__xnor2_1 _07429_ (.A(_01685_),
    .B(_01686_),
    .Y(_01689_));
 sky130_fd_sc_hd__a21o_1 _07430_ (.A1(_01688_),
    .A2(_01689_),
    .B1(_01687_),
    .X(_01690_));
 sky130_fd_sc_hd__xnor2_1 _07431_ (.A(_01681_),
    .B(_01682_),
    .Y(_01691_));
 sky130_fd_sc_hd__a21o_1 _07432_ (.A1(_01690_),
    .A2(_01691_),
    .B1(_01683_),
    .X(_01692_));
 sky130_fd_sc_hd__xnor2_1 _07433_ (.A(_01678_),
    .B(_01679_),
    .Y(_01693_));
 sky130_fd_sc_hd__a21oi_1 _07434_ (.A1(_01692_),
    .A2(_01693_),
    .B1(_01680_),
    .Y(_01694_));
 sky130_fd_sc_hd__a21o_1 _07435_ (.A1(net59),
    .A2(net25),
    .B1(_01671_),
    .X(_01696_));
 sky130_fd_sc_hd__a21boi_1 _07436_ (.A1(net59),
    .A2(_01671_),
    .B1_N(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__o311ai_1 _07437_ (.A1(_01675_),
    .A2(_01677_),
    .A3(_01697_),
    .B1(net24),
    .C1(net60),
    .Y(_01698_));
 sky130_fd_sc_hd__a2111o_1 _07438_ (.A1(net60),
    .A2(net24),
    .B1(_01675_),
    .C1(_01677_),
    .D1(_01697_),
    .X(_01699_));
 sky130_fd_sc_hd__and2_1 _07439_ (.A(_01698_),
    .B(_01699_),
    .X(_01700_));
 sky130_fd_sc_hd__nand2b_1 _07440_ (.A_N(_01694_),
    .B(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__xnor2_1 _07441_ (.A(_01694_),
    .B(_01700_),
    .Y(_01702_));
 sky130_fd_sc_hd__nand2_1 _07442_ (.A(net61),
    .B(net22),
    .Y(_01703_));
 sky130_fd_sc_hd__and3_1 _07443_ (.A(net61),
    .B(net22),
    .C(_01702_),
    .X(_01704_));
 sky130_fd_sc_hd__xor2_1 _07444_ (.A(_01692_),
    .B(_01693_),
    .X(_01705_));
 sky130_fd_sc_hd__nand2_1 _07445_ (.A(net61),
    .B(net21),
    .Y(_01707_));
 sky130_fd_sc_hd__and3_1 _07446_ (.A(net61),
    .B(net21),
    .C(_01705_),
    .X(_01708_));
 sky130_fd_sc_hd__xor2_1 _07447_ (.A(_01690_),
    .B(_01691_),
    .X(_01709_));
 sky130_fd_sc_hd__nand2_1 _07448_ (.A(net61),
    .B(net20),
    .Y(_01710_));
 sky130_fd_sc_hd__and3_1 _07449_ (.A(net61),
    .B(net20),
    .C(_01709_),
    .X(_01711_));
 sky130_fd_sc_hd__xor2_1 _07450_ (.A(_01688_),
    .B(_01689_),
    .X(_01712_));
 sky130_fd_sc_hd__nand2_1 _07451_ (.A(net61),
    .B(net19),
    .Y(_01713_));
 sky130_fd_sc_hd__and3_1 _07452_ (.A(net61),
    .B(net19),
    .C(_01712_),
    .X(_01714_));
 sky130_fd_sc_hd__a21o_1 _07453_ (.A1(_01521_),
    .A2(_01552_),
    .B1(_01551_),
    .X(_01715_));
 sky130_fd_sc_hd__xnor2_1 _07454_ (.A(_01712_),
    .B(_01713_),
    .Y(_01716_));
 sky130_fd_sc_hd__a21o_1 _07455_ (.A1(_01715_),
    .A2(_01716_),
    .B1(_01714_),
    .X(_01718_));
 sky130_fd_sc_hd__xnor2_1 _07456_ (.A(_01709_),
    .B(_01710_),
    .Y(_01719_));
 sky130_fd_sc_hd__a21o_1 _07457_ (.A1(_01718_),
    .A2(_01719_),
    .B1(_01711_),
    .X(_01720_));
 sky130_fd_sc_hd__xnor2_1 _07458_ (.A(_01705_),
    .B(_01707_),
    .Y(_01721_));
 sky130_fd_sc_hd__a21o_1 _07459_ (.A1(_01720_),
    .A2(_01721_),
    .B1(_01708_),
    .X(_01722_));
 sky130_fd_sc_hd__xnor2_1 _07460_ (.A(_01702_),
    .B(_01703_),
    .Y(_01723_));
 sky130_fd_sc_hd__a21oi_1 _07461_ (.A1(_01722_),
    .A2(_01723_),
    .B1(_01704_),
    .Y(_01724_));
 sky130_fd_sc_hd__nand2_1 _07462_ (.A(net61),
    .B(net24),
    .Y(_01725_));
 sky130_fd_sc_hd__a21o_1 _07463_ (.A1(net60),
    .A2(net25),
    .B1(_01696_),
    .X(_01726_));
 sky130_fd_sc_hd__a21bo_1 _07464_ (.A1(net60),
    .A2(_01696_),
    .B1_N(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__and3_1 _07465_ (.A(_01698_),
    .B(_01701_),
    .C(_01727_),
    .X(_01729_));
 sky130_fd_sc_hd__xnor2_1 _07466_ (.A(_01725_),
    .B(_01729_),
    .Y(_01730_));
 sky130_fd_sc_hd__or2_1 _07467_ (.A(_01724_),
    .B(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__xnor2_1 _07468_ (.A(_01724_),
    .B(_01730_),
    .Y(_01732_));
 sky130_fd_sc_hd__nand2_1 _07469_ (.A(net62),
    .B(net22),
    .Y(_01733_));
 sky130_fd_sc_hd__nor2_1 _07470_ (.A(_01732_),
    .B(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__xnor2_1 _07471_ (.A(_01722_),
    .B(_01723_),
    .Y(_01735_));
 sky130_fd_sc_hd__nand2_1 _07472_ (.A(net62),
    .B(net21),
    .Y(_01736_));
 sky130_fd_sc_hd__nor2_1 _07473_ (.A(_01735_),
    .B(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__xnor2_1 _07474_ (.A(_01720_),
    .B(_01721_),
    .Y(_01738_));
 sky130_fd_sc_hd__nand2_1 _07475_ (.A(net62),
    .B(net20),
    .Y(_01740_));
 sky130_fd_sc_hd__nor2_1 _07476_ (.A(_01738_),
    .B(_01740_),
    .Y(_01741_));
 sky130_fd_sc_hd__xnor2_1 _07477_ (.A(_01718_),
    .B(_01719_),
    .Y(_01742_));
 sky130_fd_sc_hd__nand2_1 _07478_ (.A(net62),
    .B(net19),
    .Y(_01743_));
 sky130_fd_sc_hd__nor2_1 _07479_ (.A(_01742_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__xnor2_1 _07480_ (.A(_01715_),
    .B(_01716_),
    .Y(_01745_));
 sky130_fd_sc_hd__nand2_1 _07481_ (.A(net62),
    .B(net18),
    .Y(_01746_));
 sky130_fd_sc_hd__nor2_1 _07482_ (.A(_01745_),
    .B(_01746_),
    .Y(_01747_));
 sky130_fd_sc_hd__a21o_1 _07483_ (.A1(_01518_),
    .A2(_01556_),
    .B1(_01555_),
    .X(_01748_));
 sky130_fd_sc_hd__xor2_1 _07484_ (.A(_01745_),
    .B(_01746_),
    .X(_01749_));
 sky130_fd_sc_hd__a21o_1 _07485_ (.A1(_01748_),
    .A2(_01749_),
    .B1(_01747_),
    .X(_01751_));
 sky130_fd_sc_hd__xor2_1 _07486_ (.A(_01742_),
    .B(_01743_),
    .X(_01752_));
 sky130_fd_sc_hd__a21o_1 _07487_ (.A1(_01751_),
    .A2(_01752_),
    .B1(_01744_),
    .X(_01753_));
 sky130_fd_sc_hd__xor2_1 _07488_ (.A(_01738_),
    .B(_01740_),
    .X(_01754_));
 sky130_fd_sc_hd__a21o_1 _07489_ (.A1(_01753_),
    .A2(_01754_),
    .B1(_01741_),
    .X(_01755_));
 sky130_fd_sc_hd__xor2_1 _07490_ (.A(_01735_),
    .B(_01736_),
    .X(_01756_));
 sky130_fd_sc_hd__a21o_1 _07491_ (.A1(_01755_),
    .A2(_01756_),
    .B1(_01737_),
    .X(_01757_));
 sky130_fd_sc_hd__xor2_1 _07492_ (.A(_01732_),
    .B(_01733_),
    .X(_01758_));
 sky130_fd_sc_hd__a21oi_1 _07493_ (.A1(_01757_),
    .A2(_01758_),
    .B1(_01734_),
    .Y(_01759_));
 sky130_fd_sc_hd__a21o_1 _07494_ (.A1(net61),
    .A2(net25),
    .B1(_01726_),
    .X(_01760_));
 sky130_fd_sc_hd__inv_2 _07495_ (.A(_01760_),
    .Y(_01762_));
 sky130_fd_sc_hd__and3_1 _07496_ (.A(net61),
    .B(net25),
    .C(_01726_),
    .X(_01763_));
 sky130_fd_sc_hd__o221a_1 _07497_ (.A1(_01725_),
    .A2(_01729_),
    .B1(_01762_),
    .B2(_01763_),
    .C1(_01731_),
    .X(_01764_));
 sky130_fd_sc_hd__nand2_1 _07498_ (.A(net62),
    .B(net24),
    .Y(_01765_));
 sky130_fd_sc_hd__xnor2_1 _07499_ (.A(_01764_),
    .B(_01765_),
    .Y(_01766_));
 sky130_fd_sc_hd__xnor2_1 _07500_ (.A(_01759_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__nand2_1 _07501_ (.A(net63),
    .B(net22),
    .Y(_01768_));
 sky130_fd_sc_hd__nor2_1 _07502_ (.A(_01767_),
    .B(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__xnor2_1 _07503_ (.A(_01757_),
    .B(_01758_),
    .Y(_01770_));
 sky130_fd_sc_hd__nand2_1 _07504_ (.A(net63),
    .B(net21),
    .Y(_01771_));
 sky130_fd_sc_hd__nor2_1 _07505_ (.A(_01770_),
    .B(_01771_),
    .Y(_01773_));
 sky130_fd_sc_hd__xnor2_1 _07506_ (.A(_01755_),
    .B(_01756_),
    .Y(_01774_));
 sky130_fd_sc_hd__nand2_1 _07507_ (.A(net63),
    .B(net20),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2_1 _07508_ (.A(_01774_),
    .B(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__xnor2_1 _07509_ (.A(_01753_),
    .B(_01754_),
    .Y(_01777_));
 sky130_fd_sc_hd__nand2_1 _07510_ (.A(net63),
    .B(net19),
    .Y(_01778_));
 sky130_fd_sc_hd__nor2_1 _07511_ (.A(_01777_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__xnor2_1 _07512_ (.A(_01751_),
    .B(_01752_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand2_1 _07513_ (.A(net63),
    .B(net18),
    .Y(_01781_));
 sky130_fd_sc_hd__nor2_1 _07514_ (.A(_01780_),
    .B(_01781_),
    .Y(_01782_));
 sky130_fd_sc_hd__xnor2_1 _07515_ (.A(_01748_),
    .B(_01749_),
    .Y(_01784_));
 sky130_fd_sc_hd__nand2_1 _07516_ (.A(net63),
    .B(net17),
    .Y(_01785_));
 sky130_fd_sc_hd__nor2_1 _07517_ (.A(_01784_),
    .B(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__a21o_1 _07518_ (.A1(_01516_),
    .A2(_01559_),
    .B1(_01558_),
    .X(_01787_));
 sky130_fd_sc_hd__xor2_1 _07519_ (.A(_01784_),
    .B(_01785_),
    .X(_01788_));
 sky130_fd_sc_hd__a21o_1 _07520_ (.A1(_01787_),
    .A2(_01788_),
    .B1(_01786_),
    .X(_01789_));
 sky130_fd_sc_hd__xor2_1 _07521_ (.A(_01780_),
    .B(_01781_),
    .X(_01790_));
 sky130_fd_sc_hd__a21o_1 _07522_ (.A1(_01789_),
    .A2(_01790_),
    .B1(_01782_),
    .X(_01791_));
 sky130_fd_sc_hd__xor2_1 _07523_ (.A(_01777_),
    .B(_01778_),
    .X(_01792_));
 sky130_fd_sc_hd__a21o_1 _07524_ (.A1(_01791_),
    .A2(_01792_),
    .B1(_01779_),
    .X(_01793_));
 sky130_fd_sc_hd__xor2_1 _07525_ (.A(_01774_),
    .B(_01775_),
    .X(_01795_));
 sky130_fd_sc_hd__a21o_1 _07526_ (.A1(_01793_),
    .A2(_01795_),
    .B1(_01776_),
    .X(_01796_));
 sky130_fd_sc_hd__xor2_1 _07527_ (.A(_01770_),
    .B(_01771_),
    .X(_01797_));
 sky130_fd_sc_hd__a21o_1 _07528_ (.A1(_01796_),
    .A2(_01797_),
    .B1(_01773_),
    .X(_01798_));
 sky130_fd_sc_hd__xor2_1 _07529_ (.A(_01767_),
    .B(_01768_),
    .X(_01799_));
 sky130_fd_sc_hd__a21oi_1 _07530_ (.A1(_01798_),
    .A2(_01799_),
    .B1(_01769_),
    .Y(_01800_));
 sky130_fd_sc_hd__nand2_1 _07531_ (.A(net62),
    .B(net25),
    .Y(_01801_));
 sky130_fd_sc_hd__and2_1 _07532_ (.A(_01762_),
    .B(_01801_),
    .X(_01802_));
 sky130_fd_sc_hd__nor2_1 _07533_ (.A(_01762_),
    .B(_01801_),
    .Y(_01803_));
 sky130_fd_sc_hd__o22a_1 _07534_ (.A1(_01759_),
    .A2(_01766_),
    .B1(_01802_),
    .B2(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__o21ai_1 _07535_ (.A1(_01764_),
    .A2(_01765_),
    .B1(_01804_),
    .Y(_01806_));
 sky130_fd_sc_hd__nand2_1 _07536_ (.A(net63),
    .B(net24),
    .Y(_01807_));
 sky130_fd_sc_hd__xor2_1 _07537_ (.A(_01806_),
    .B(_01807_),
    .X(_01808_));
 sky130_fd_sc_hd__xnor2_1 _07538_ (.A(_01800_),
    .B(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__nand2_1 _07539_ (.A(net64),
    .B(net22),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_1 _07540_ (.A(_01809_),
    .B(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__xnor2_1 _07541_ (.A(_01798_),
    .B(_01799_),
    .Y(_01812_));
 sky130_fd_sc_hd__nand2_1 _07542_ (.A(net64),
    .B(net21),
    .Y(_01813_));
 sky130_fd_sc_hd__nor2_1 _07543_ (.A(_01812_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__xnor2_1 _07544_ (.A(_01796_),
    .B(_01797_),
    .Y(_01815_));
 sky130_fd_sc_hd__nand2_1 _07545_ (.A(net64),
    .B(net20),
    .Y(_01817_));
 sky130_fd_sc_hd__nor2_1 _07546_ (.A(_01815_),
    .B(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__xnor2_1 _07547_ (.A(_01793_),
    .B(_01795_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand2_1 _07548_ (.A(net64),
    .B(net19),
    .Y(_01820_));
 sky130_fd_sc_hd__nor2_1 _07549_ (.A(_01819_),
    .B(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__xnor2_1 _07550_ (.A(_01791_),
    .B(_01792_),
    .Y(_01822_));
 sky130_fd_sc_hd__nand2_1 _07551_ (.A(net64),
    .B(net18),
    .Y(_01823_));
 sky130_fd_sc_hd__nor2_1 _07552_ (.A(_01822_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__xnor2_1 _07553_ (.A(_01789_),
    .B(_01790_),
    .Y(_01825_));
 sky130_fd_sc_hd__nand2_1 _07554_ (.A(net64),
    .B(net17),
    .Y(_01826_));
 sky130_fd_sc_hd__nor2_1 _07555_ (.A(_01825_),
    .B(_01826_),
    .Y(_01828_));
 sky130_fd_sc_hd__xnor2_1 _07556_ (.A(_01787_),
    .B(_01788_),
    .Y(_01829_));
 sky130_fd_sc_hd__nand2_1 _07557_ (.A(net64),
    .B(net16),
    .Y(_01830_));
 sky130_fd_sc_hd__nor2_1 _07558_ (.A(_01829_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__a21o_1 _07559_ (.A1(_01514_),
    .A2(_01562_),
    .B1(_01561_),
    .X(_01832_));
 sky130_fd_sc_hd__xor2_1 _07560_ (.A(_01829_),
    .B(_01830_),
    .X(_01833_));
 sky130_fd_sc_hd__a21o_1 _07561_ (.A1(_01832_),
    .A2(_01833_),
    .B1(_01831_),
    .X(_01834_));
 sky130_fd_sc_hd__xor2_1 _07562_ (.A(_01825_),
    .B(_01826_),
    .X(_01835_));
 sky130_fd_sc_hd__a21o_1 _07563_ (.A1(_01834_),
    .A2(_01835_),
    .B1(_01828_),
    .X(_01836_));
 sky130_fd_sc_hd__xor2_1 _07564_ (.A(_01822_),
    .B(_01823_),
    .X(_01837_));
 sky130_fd_sc_hd__a21o_1 _07565_ (.A1(_01836_),
    .A2(_01837_),
    .B1(_01824_),
    .X(_01839_));
 sky130_fd_sc_hd__xor2_1 _07566_ (.A(_01819_),
    .B(_01820_),
    .X(_01840_));
 sky130_fd_sc_hd__a21o_1 _07567_ (.A1(_01839_),
    .A2(_01840_),
    .B1(_01821_),
    .X(_01841_));
 sky130_fd_sc_hd__xor2_1 _07568_ (.A(_01815_),
    .B(_01817_),
    .X(_01842_));
 sky130_fd_sc_hd__a21o_1 _07569_ (.A1(_01841_),
    .A2(_01842_),
    .B1(_01818_),
    .X(_01843_));
 sky130_fd_sc_hd__xor2_1 _07570_ (.A(_01812_),
    .B(_01813_),
    .X(_01844_));
 sky130_fd_sc_hd__a21o_1 _07571_ (.A1(_01843_),
    .A2(_01844_),
    .B1(_01814_),
    .X(_01845_));
 sky130_fd_sc_hd__xor2_1 _07572_ (.A(_01809_),
    .B(_01810_),
    .X(_01846_));
 sky130_fd_sc_hd__a21oi_1 _07573_ (.A1(_01845_),
    .A2(_01846_),
    .B1(_01811_),
    .Y(_01847_));
 sky130_fd_sc_hd__nand2_1 _07574_ (.A(net63),
    .B(net25),
    .Y(_01848_));
 sky130_fd_sc_hd__nand2_1 _07575_ (.A(_01802_),
    .B(_01848_),
    .Y(_01850_));
 sky130_fd_sc_hd__or2_1 _07576_ (.A(_01802_),
    .B(_01848_),
    .X(_01851_));
 sky130_fd_sc_hd__a2bb2o_1 _07577_ (.A1_N(_01800_),
    .A2_N(_01808_),
    .B1(_01850_),
    .B2(_01851_),
    .X(_01852_));
 sky130_fd_sc_hd__a31o_1 _07578_ (.A1(net63),
    .A2(net24),
    .A3(_01806_),
    .B1(_01852_),
    .X(_01853_));
 sky130_fd_sc_hd__nand2_1 _07579_ (.A(net64),
    .B(net24),
    .Y(_01854_));
 sky130_fd_sc_hd__and3_1 _07580_ (.A(net64),
    .B(net24),
    .C(_01853_),
    .X(_01855_));
 sky130_fd_sc_hd__xor2_1 _07581_ (.A(_01853_),
    .B(_01854_),
    .X(_01856_));
 sky130_fd_sc_hd__xnor2_1 _07582_ (.A(_01847_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__nand2_1 _07583_ (.A(net34),
    .B(net22),
    .Y(_01858_));
 sky130_fd_sc_hd__nor2_1 _07584_ (.A(_01857_),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__xnor2_1 _07585_ (.A(_01845_),
    .B(_01846_),
    .Y(_01861_));
 sky130_fd_sc_hd__nand2_1 _07586_ (.A(net34),
    .B(net21),
    .Y(_01862_));
 sky130_fd_sc_hd__nor2_1 _07587_ (.A(_01861_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__xnor2_1 _07588_ (.A(_01843_),
    .B(_01844_),
    .Y(_01864_));
 sky130_fd_sc_hd__nand2_1 _07589_ (.A(net34),
    .B(net20),
    .Y(_01865_));
 sky130_fd_sc_hd__nor2_1 _07590_ (.A(_01864_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__xnor2_1 _07591_ (.A(_01841_),
    .B(_01842_),
    .Y(_01867_));
 sky130_fd_sc_hd__nand2_1 _07592_ (.A(net34),
    .B(net19),
    .Y(_01868_));
 sky130_fd_sc_hd__nor2_1 _07593_ (.A(_01867_),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__xnor2_1 _07594_ (.A(_01839_),
    .B(_01840_),
    .Y(_01870_));
 sky130_fd_sc_hd__nand2_1 _07595_ (.A(net34),
    .B(net18),
    .Y(_01872_));
 sky130_fd_sc_hd__nor2_1 _07596_ (.A(_01870_),
    .B(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__xnor2_1 _07597_ (.A(_01836_),
    .B(_01837_),
    .Y(_01874_));
 sky130_fd_sc_hd__nand2_1 _07598_ (.A(net34),
    .B(net17),
    .Y(_01875_));
 sky130_fd_sc_hd__nor2_1 _07599_ (.A(_01874_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__xnor2_1 _07600_ (.A(_01834_),
    .B(_01835_),
    .Y(_01877_));
 sky130_fd_sc_hd__nand2_1 _07601_ (.A(net34),
    .B(net16),
    .Y(_01878_));
 sky130_fd_sc_hd__nor2_1 _07602_ (.A(_01877_),
    .B(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__xnor2_1 _07603_ (.A(_01832_),
    .B(_01833_),
    .Y(_01880_));
 sky130_fd_sc_hd__nand2_1 _07604_ (.A(net34),
    .B(net15),
    .Y(_01881_));
 sky130_fd_sc_hd__nor2_1 _07605_ (.A(_01880_),
    .B(_01881_),
    .Y(_01883_));
 sky130_fd_sc_hd__a21o_1 _07606_ (.A1(_01512_),
    .A2(_01566_),
    .B1(_01565_),
    .X(_01884_));
 sky130_fd_sc_hd__xor2_1 _07607_ (.A(_01880_),
    .B(_01881_),
    .X(_01885_));
 sky130_fd_sc_hd__a21o_1 _07608_ (.A1(_01884_),
    .A2(_01885_),
    .B1(_01883_),
    .X(_01886_));
 sky130_fd_sc_hd__xor2_1 _07609_ (.A(_01877_),
    .B(_01878_),
    .X(_01887_));
 sky130_fd_sc_hd__a21o_1 _07610_ (.A1(_01886_),
    .A2(_01887_),
    .B1(_01879_),
    .X(_01888_));
 sky130_fd_sc_hd__xor2_1 _07611_ (.A(_01874_),
    .B(_01875_),
    .X(_01889_));
 sky130_fd_sc_hd__a21o_1 _07612_ (.A1(_01888_),
    .A2(_01889_),
    .B1(_01876_),
    .X(_01890_));
 sky130_fd_sc_hd__xor2_1 _07613_ (.A(_01870_),
    .B(_01872_),
    .X(_01891_));
 sky130_fd_sc_hd__a21o_1 _07614_ (.A1(_01890_),
    .A2(_01891_),
    .B1(_01873_),
    .X(_01892_));
 sky130_fd_sc_hd__xor2_1 _07615_ (.A(_01867_),
    .B(_01868_),
    .X(_01894_));
 sky130_fd_sc_hd__a21o_1 _07616_ (.A1(_01892_),
    .A2(_01894_),
    .B1(_01869_),
    .X(_01895_));
 sky130_fd_sc_hd__xor2_1 _07617_ (.A(_01864_),
    .B(_01865_),
    .X(_01896_));
 sky130_fd_sc_hd__a21o_1 _07618_ (.A1(_01895_),
    .A2(_01896_),
    .B1(_01866_),
    .X(_01897_));
 sky130_fd_sc_hd__xor2_1 _07619_ (.A(_01861_),
    .B(_01862_),
    .X(_01898_));
 sky130_fd_sc_hd__a21o_1 _07620_ (.A1(_01897_),
    .A2(_01898_),
    .B1(_01863_),
    .X(_01899_));
 sky130_fd_sc_hd__xor2_1 _07621_ (.A(_01857_),
    .B(_01858_),
    .X(_01900_));
 sky130_fd_sc_hd__a21oi_1 _07622_ (.A1(_01899_),
    .A2(_01900_),
    .B1(_01859_),
    .Y(_01901_));
 sky130_fd_sc_hd__nand2_1 _07623_ (.A(net64),
    .B(net25),
    .Y(_01902_));
 sky130_fd_sc_hd__and3_1 _07624_ (.A(_01802_),
    .B(_01848_),
    .C(_01902_),
    .X(_01903_));
 sky130_fd_sc_hd__and3_1 _07625_ (.A(net64),
    .B(net25),
    .C(_01850_),
    .X(_01905_));
 sky130_fd_sc_hd__o21ba_1 _07626_ (.A1(_01847_),
    .A2(_01856_),
    .B1_N(_01855_),
    .X(_01906_));
 sky130_fd_sc_hd__o21ai_1 _07627_ (.A1(_01903_),
    .A2(_01905_),
    .B1(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _07628_ (.A(net34),
    .B(net24),
    .Y(_01908_));
 sky130_fd_sc_hd__and3_1 _07629_ (.A(net34),
    .B(net24),
    .C(_01907_),
    .X(_01909_));
 sky130_fd_sc_hd__xor2_1 _07630_ (.A(_01907_),
    .B(_01908_),
    .X(_01910_));
 sky130_fd_sc_hd__xnor2_1 _07631_ (.A(_01901_),
    .B(_01910_),
    .Y(_01911_));
 sky130_fd_sc_hd__nand2_1 _07632_ (.A(net35),
    .B(net22),
    .Y(_01912_));
 sky130_fd_sc_hd__nor2_1 _07633_ (.A(_01911_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__xnor2_1 _07634_ (.A(_01899_),
    .B(_01900_),
    .Y(_01914_));
 sky130_fd_sc_hd__nand2_1 _07635_ (.A(net35),
    .B(net21),
    .Y(_01916_));
 sky130_fd_sc_hd__nor2_1 _07636_ (.A(_01914_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__xnor2_1 _07637_ (.A(_01897_),
    .B(_01898_),
    .Y(_01918_));
 sky130_fd_sc_hd__nand2_1 _07638_ (.A(net35),
    .B(net20),
    .Y(_01919_));
 sky130_fd_sc_hd__nor2_1 _07639_ (.A(_01918_),
    .B(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hd__xnor2_1 _07640_ (.A(_01895_),
    .B(_01896_),
    .Y(_01921_));
 sky130_fd_sc_hd__nand2_1 _07641_ (.A(net35),
    .B(net19),
    .Y(_01922_));
 sky130_fd_sc_hd__nor2_1 _07642_ (.A(_01921_),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__xnor2_1 _07643_ (.A(_01892_),
    .B(_01894_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand2_1 _07644_ (.A(net35),
    .B(net18),
    .Y(_01925_));
 sky130_fd_sc_hd__nor2_1 _07645_ (.A(_01924_),
    .B(_01925_),
    .Y(_01927_));
 sky130_fd_sc_hd__xnor2_1 _07646_ (.A(_01890_),
    .B(_01891_),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_1 _07647_ (.A(net35),
    .B(net17),
    .Y(_01929_));
 sky130_fd_sc_hd__nor2_1 _07648_ (.A(_01928_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__xnor2_1 _07649_ (.A(_01888_),
    .B(_01889_),
    .Y(_01931_));
 sky130_fd_sc_hd__nand2_1 _07650_ (.A(net35),
    .B(net16),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_1 _07651_ (.A(_01931_),
    .B(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__xnor2_1 _07652_ (.A(_01886_),
    .B(_01887_),
    .Y(_01934_));
 sky130_fd_sc_hd__nand2_1 _07653_ (.A(net35),
    .B(net15),
    .Y(_01935_));
 sky130_fd_sc_hd__nor2_1 _07654_ (.A(_01934_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__xnor2_1 _07655_ (.A(_01884_),
    .B(_01885_),
    .Y(_01938_));
 sky130_fd_sc_hd__nand2_1 _07656_ (.A(net35),
    .B(net14),
    .Y(_01939_));
 sky130_fd_sc_hd__nor2_1 _07657_ (.A(_01938_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__a21o_1 _07658_ (.A1(_01510_),
    .A2(_01569_),
    .B1(_01568_),
    .X(_01941_));
 sky130_fd_sc_hd__xor2_1 _07659_ (.A(_01938_),
    .B(_01939_),
    .X(_01942_));
 sky130_fd_sc_hd__a21o_1 _07660_ (.A1(_01941_),
    .A2(_01942_),
    .B1(_01940_),
    .X(_01943_));
 sky130_fd_sc_hd__xor2_1 _07661_ (.A(_01934_),
    .B(_01935_),
    .X(_01944_));
 sky130_fd_sc_hd__a21o_1 _07662_ (.A1(_01943_),
    .A2(_01944_),
    .B1(_01936_),
    .X(_01945_));
 sky130_fd_sc_hd__xor2_1 _07663_ (.A(_01931_),
    .B(_01932_),
    .X(_01946_));
 sky130_fd_sc_hd__a21o_1 _07664_ (.A1(_01945_),
    .A2(_01946_),
    .B1(_01933_),
    .X(_01947_));
 sky130_fd_sc_hd__xor2_1 _07665_ (.A(_01928_),
    .B(_01929_),
    .X(_01949_));
 sky130_fd_sc_hd__a21o_1 _07666_ (.A1(_01947_),
    .A2(_01949_),
    .B1(_01930_),
    .X(_01950_));
 sky130_fd_sc_hd__xor2_1 _07667_ (.A(_01924_),
    .B(_01925_),
    .X(_01951_));
 sky130_fd_sc_hd__a21o_1 _07668_ (.A1(_01950_),
    .A2(_01951_),
    .B1(_01927_),
    .X(_01952_));
 sky130_fd_sc_hd__xor2_1 _07669_ (.A(_01921_),
    .B(_01922_),
    .X(_01953_));
 sky130_fd_sc_hd__a21o_1 _07670_ (.A1(_01952_),
    .A2(_01953_),
    .B1(_01923_),
    .X(_01954_));
 sky130_fd_sc_hd__xor2_1 _07671_ (.A(_01918_),
    .B(_01919_),
    .X(_01955_));
 sky130_fd_sc_hd__a21o_1 _07672_ (.A1(_01954_),
    .A2(_01955_),
    .B1(_01920_),
    .X(_01956_));
 sky130_fd_sc_hd__xor2_1 _07673_ (.A(_01914_),
    .B(_01916_),
    .X(_01957_));
 sky130_fd_sc_hd__a21o_1 _07674_ (.A1(_01956_),
    .A2(_01957_),
    .B1(_01917_),
    .X(_01958_));
 sky130_fd_sc_hd__xor2_1 _07675_ (.A(_01911_),
    .B(_01912_),
    .X(_01960_));
 sky130_fd_sc_hd__a21oi_1 _07676_ (.A1(_01958_),
    .A2(_01960_),
    .B1(_01913_),
    .Y(_01961_));
 sky130_fd_sc_hd__nand2_1 _07677_ (.A(net34),
    .B(net25),
    .Y(_01962_));
 sky130_fd_sc_hd__and2_1 _07678_ (.A(_01903_),
    .B(_01962_),
    .X(_01963_));
 sky130_fd_sc_hd__nor2_1 _07679_ (.A(_01903_),
    .B(_01962_),
    .Y(_01964_));
 sky130_fd_sc_hd__o21ba_1 _07680_ (.A1(_01901_),
    .A2(_01910_),
    .B1_N(_01909_),
    .X(_01965_));
 sky130_fd_sc_hd__o21ai_1 _07681_ (.A1(_01963_),
    .A2(_01964_),
    .B1(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__nand2_1 _07682_ (.A(net35),
    .B(net24),
    .Y(_01967_));
 sky130_fd_sc_hd__xor2_1 _07683_ (.A(_01966_),
    .B(_01967_),
    .X(_01968_));
 sky130_fd_sc_hd__xnor2_1 _07684_ (.A(_01961_),
    .B(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__nand2_1 _07685_ (.A(net36),
    .B(net22),
    .Y(_01971_));
 sky130_fd_sc_hd__nor2_1 _07686_ (.A(_01969_),
    .B(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__xnor2_1 _07687_ (.A(_01958_),
    .B(_01960_),
    .Y(_01973_));
 sky130_fd_sc_hd__nand2_1 _07688_ (.A(net36),
    .B(net21),
    .Y(_01974_));
 sky130_fd_sc_hd__nor2_1 _07689_ (.A(_01973_),
    .B(_01974_),
    .Y(_01975_));
 sky130_fd_sc_hd__xnor2_1 _07690_ (.A(_01956_),
    .B(_01957_),
    .Y(_01976_));
 sky130_fd_sc_hd__nand2_1 _07691_ (.A(net36),
    .B(net20),
    .Y(_01977_));
 sky130_fd_sc_hd__nor2_1 _07692_ (.A(_01976_),
    .B(_01977_),
    .Y(_01978_));
 sky130_fd_sc_hd__xnor2_1 _07693_ (.A(_01954_),
    .B(_01955_),
    .Y(_01979_));
 sky130_fd_sc_hd__nand2_1 _07694_ (.A(net36),
    .B(net19),
    .Y(_01980_));
 sky130_fd_sc_hd__nor2_1 _07695_ (.A(_01979_),
    .B(_01980_),
    .Y(_01982_));
 sky130_fd_sc_hd__xnor2_1 _07696_ (.A(_01952_),
    .B(_01953_),
    .Y(_01983_));
 sky130_fd_sc_hd__nand2_1 _07697_ (.A(net36),
    .B(net18),
    .Y(_01984_));
 sky130_fd_sc_hd__nor2_1 _07698_ (.A(_01983_),
    .B(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__xnor2_1 _07699_ (.A(_01950_),
    .B(_01951_),
    .Y(_01986_));
 sky130_fd_sc_hd__nand2_1 _07700_ (.A(net36),
    .B(net17),
    .Y(_01987_));
 sky130_fd_sc_hd__nor2_1 _07701_ (.A(_01986_),
    .B(_01987_),
    .Y(_01988_));
 sky130_fd_sc_hd__xnor2_1 _07702_ (.A(_01947_),
    .B(_01949_),
    .Y(_01989_));
 sky130_fd_sc_hd__nand2_1 _07703_ (.A(net36),
    .B(net16),
    .Y(_01990_));
 sky130_fd_sc_hd__nor2_1 _07704_ (.A(_01989_),
    .B(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__xnor2_1 _07705_ (.A(_01945_),
    .B(_01946_),
    .Y(_01993_));
 sky130_fd_sc_hd__nand2_1 _07706_ (.A(net36),
    .B(net15),
    .Y(_01994_));
 sky130_fd_sc_hd__nor2_1 _07707_ (.A(_01993_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__xnor2_1 _07708_ (.A(_01943_),
    .B(_01944_),
    .Y(_01996_));
 sky130_fd_sc_hd__nand2_1 _07709_ (.A(net36),
    .B(net14),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_1 _07710_ (.A(_01996_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__xnor2_1 _07711_ (.A(_01941_),
    .B(_01942_),
    .Y(_01999_));
 sky130_fd_sc_hd__nand2_1 _07712_ (.A(net36),
    .B(net13),
    .Y(_02000_));
 sky130_fd_sc_hd__nor2_1 _07713_ (.A(_01999_),
    .B(_02000_),
    .Y(_02001_));
 sky130_fd_sc_hd__a21o_1 _07714_ (.A1(_01507_),
    .A2(_01572_),
    .B1(_01571_),
    .X(_02002_));
 sky130_fd_sc_hd__xor2_1 _07715_ (.A(_01999_),
    .B(_02000_),
    .X(_02004_));
 sky130_fd_sc_hd__a21o_1 _07716_ (.A1(_02002_),
    .A2(_02004_),
    .B1(_02001_),
    .X(_02005_));
 sky130_fd_sc_hd__xor2_1 _07717_ (.A(_01996_),
    .B(_01997_),
    .X(_02006_));
 sky130_fd_sc_hd__a21o_1 _07718_ (.A1(_02005_),
    .A2(_02006_),
    .B1(_01998_),
    .X(_02007_));
 sky130_fd_sc_hd__xor2_1 _07719_ (.A(_01993_),
    .B(_01994_),
    .X(_02008_));
 sky130_fd_sc_hd__a21o_1 _07720_ (.A1(_02007_),
    .A2(_02008_),
    .B1(_01995_),
    .X(_02009_));
 sky130_fd_sc_hd__xor2_1 _07721_ (.A(_01989_),
    .B(_01990_),
    .X(_02010_));
 sky130_fd_sc_hd__a21o_1 _07722_ (.A1(_02009_),
    .A2(_02010_),
    .B1(_01991_),
    .X(_02011_));
 sky130_fd_sc_hd__xor2_1 _07723_ (.A(_01986_),
    .B(_01987_),
    .X(_02012_));
 sky130_fd_sc_hd__a21o_1 _07724_ (.A1(_02011_),
    .A2(_02012_),
    .B1(_01988_),
    .X(_02013_));
 sky130_fd_sc_hd__xor2_1 _07725_ (.A(_01983_),
    .B(_01984_),
    .X(_02015_));
 sky130_fd_sc_hd__a21o_1 _07726_ (.A1(_02013_),
    .A2(_02015_),
    .B1(_01985_),
    .X(_02016_));
 sky130_fd_sc_hd__xor2_1 _07727_ (.A(_01979_),
    .B(_01980_),
    .X(_02017_));
 sky130_fd_sc_hd__a21o_1 _07728_ (.A1(_02016_),
    .A2(_02017_),
    .B1(_01982_),
    .X(_02018_));
 sky130_fd_sc_hd__xor2_1 _07729_ (.A(_01976_),
    .B(_01977_),
    .X(_02019_));
 sky130_fd_sc_hd__a21o_1 _07730_ (.A1(_02018_),
    .A2(_02019_),
    .B1(_01978_),
    .X(_02020_));
 sky130_fd_sc_hd__xor2_1 _07731_ (.A(_01973_),
    .B(_01974_),
    .X(_02021_));
 sky130_fd_sc_hd__a21o_1 _07732_ (.A1(_02020_),
    .A2(_02021_),
    .B1(_01975_),
    .X(_02022_));
 sky130_fd_sc_hd__xor2_1 _07733_ (.A(_01969_),
    .B(_01971_),
    .X(_02023_));
 sky130_fd_sc_hd__a21oi_1 _07734_ (.A1(_02022_),
    .A2(_02023_),
    .B1(_01972_),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_1 _07735_ (.A(net35),
    .B(net25),
    .Y(_02026_));
 sky130_fd_sc_hd__nand2_1 _07736_ (.A(_01963_),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__or2_1 _07737_ (.A(_01963_),
    .B(_02026_),
    .X(_02028_));
 sky130_fd_sc_hd__a2bb2o_1 _07738_ (.A1_N(_01961_),
    .A2_N(_01968_),
    .B1(_02027_),
    .B2(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__a31o_1 _07739_ (.A1(net35),
    .A2(net24),
    .A3(_01966_),
    .B1(_02029_),
    .X(_02030_));
 sky130_fd_sc_hd__nand2_1 _07740_ (.A(net36),
    .B(net24),
    .Y(_02031_));
 sky130_fd_sc_hd__and3_1 _07741_ (.A(net36),
    .B(net24),
    .C(_02030_),
    .X(_02032_));
 sky130_fd_sc_hd__xor2_1 _07742_ (.A(_02030_),
    .B(_02031_),
    .X(_02033_));
 sky130_fd_sc_hd__xnor2_1 _07743_ (.A(_02024_),
    .B(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _07744_ (.A(net37),
    .B(net22),
    .Y(_02035_));
 sky130_fd_sc_hd__nor2_1 _07745_ (.A(_02034_),
    .B(_02035_),
    .Y(_02037_));
 sky130_fd_sc_hd__xnor2_1 _07746_ (.A(_02022_),
    .B(_02023_),
    .Y(_02038_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(net37),
    .B(net21),
    .Y(_02039_));
 sky130_fd_sc_hd__nor2_1 _07748_ (.A(_02038_),
    .B(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__xnor2_1 _07749_ (.A(_02020_),
    .B(_02021_),
    .Y(_02041_));
 sky130_fd_sc_hd__nand2_1 _07750_ (.A(net37),
    .B(net20),
    .Y(_02042_));
 sky130_fd_sc_hd__nor2_1 _07751_ (.A(_02041_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__xnor2_1 _07752_ (.A(_02018_),
    .B(_02019_),
    .Y(_02044_));
 sky130_fd_sc_hd__nand2_1 _07753_ (.A(net37),
    .B(net19),
    .Y(_02045_));
 sky130_fd_sc_hd__nor2_1 _07754_ (.A(_02044_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__xnor2_1 _07755_ (.A(_02016_),
    .B(_02017_),
    .Y(_02048_));
 sky130_fd_sc_hd__nand2_1 _07756_ (.A(net37),
    .B(net18),
    .Y(_02049_));
 sky130_fd_sc_hd__nor2_1 _07757_ (.A(_02048_),
    .B(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__xnor2_1 _07758_ (.A(_02013_),
    .B(_02015_),
    .Y(_02051_));
 sky130_fd_sc_hd__nand2_1 _07759_ (.A(net37),
    .B(net17),
    .Y(_02052_));
 sky130_fd_sc_hd__nor2_1 _07760_ (.A(_02051_),
    .B(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__xnor2_1 _07761_ (.A(_02011_),
    .B(_02012_),
    .Y(_02054_));
 sky130_fd_sc_hd__nand2_1 _07762_ (.A(net37),
    .B(net16),
    .Y(_02055_));
 sky130_fd_sc_hd__nor2_1 _07763_ (.A(_02054_),
    .B(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__xnor2_1 _07764_ (.A(_02009_),
    .B(_02010_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2_1 _07765_ (.A(net37),
    .B(net15),
    .Y(_02059_));
 sky130_fd_sc_hd__nor2_1 _07766_ (.A(_02057_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__xnor2_1 _07767_ (.A(_02007_),
    .B(_02008_),
    .Y(_02061_));
 sky130_fd_sc_hd__nand2_1 _07768_ (.A(net37),
    .B(net14),
    .Y(_02062_));
 sky130_fd_sc_hd__nor2_1 _07769_ (.A(_02061_),
    .B(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__xnor2_1 _07770_ (.A(_02005_),
    .B(_02006_),
    .Y(_02064_));
 sky130_fd_sc_hd__nand2_1 _07771_ (.A(net37),
    .B(net13),
    .Y(_02065_));
 sky130_fd_sc_hd__nor2_1 _07772_ (.A(_02064_),
    .B(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__xnor2_1 _07773_ (.A(_02002_),
    .B(_02004_),
    .Y(_02067_));
 sky130_fd_sc_hd__nand2_1 _07774_ (.A(net37),
    .B(net11),
    .Y(_02068_));
 sky130_fd_sc_hd__nor2_1 _07775_ (.A(_02067_),
    .B(_02068_),
    .Y(_02070_));
 sky130_fd_sc_hd__a21o_1 _07776_ (.A1(_01505_),
    .A2(_01576_),
    .B1(_01574_),
    .X(_02071_));
 sky130_fd_sc_hd__xor2_1 _07777_ (.A(_02067_),
    .B(_02068_),
    .X(_02072_));
 sky130_fd_sc_hd__a21o_1 _07778_ (.A1(_02071_),
    .A2(_02072_),
    .B1(_02070_),
    .X(_02073_));
 sky130_fd_sc_hd__xor2_1 _07779_ (.A(_02064_),
    .B(_02065_),
    .X(_02074_));
 sky130_fd_sc_hd__a21o_1 _07780_ (.A1(_02073_),
    .A2(_02074_),
    .B1(_02066_),
    .X(_02075_));
 sky130_fd_sc_hd__xor2_1 _07781_ (.A(_02061_),
    .B(_02062_),
    .X(_02076_));
 sky130_fd_sc_hd__a21o_1 _07782_ (.A1(_02075_),
    .A2(_02076_),
    .B1(_02063_),
    .X(_02077_));
 sky130_fd_sc_hd__xor2_1 _07783_ (.A(_02057_),
    .B(_02059_),
    .X(_02078_));
 sky130_fd_sc_hd__a21o_1 _07784_ (.A1(_02077_),
    .A2(_02078_),
    .B1(_02060_),
    .X(_02079_));
 sky130_fd_sc_hd__xor2_1 _07785_ (.A(_02054_),
    .B(_02055_),
    .X(_02081_));
 sky130_fd_sc_hd__a21o_1 _07786_ (.A1(_02079_),
    .A2(_02081_),
    .B1(_02056_),
    .X(_02082_));
 sky130_fd_sc_hd__xor2_1 _07787_ (.A(_02051_),
    .B(_02052_),
    .X(_02083_));
 sky130_fd_sc_hd__a21o_1 _07788_ (.A1(_02082_),
    .A2(_02083_),
    .B1(_02053_),
    .X(_02084_));
 sky130_fd_sc_hd__xor2_1 _07789_ (.A(_02048_),
    .B(_02049_),
    .X(_02085_));
 sky130_fd_sc_hd__a21o_1 _07790_ (.A1(_02084_),
    .A2(_02085_),
    .B1(_02050_),
    .X(_02086_));
 sky130_fd_sc_hd__xor2_1 _07791_ (.A(_02044_),
    .B(_02045_),
    .X(_02087_));
 sky130_fd_sc_hd__a21o_1 _07792_ (.A1(_02086_),
    .A2(_02087_),
    .B1(_02046_),
    .X(_02088_));
 sky130_fd_sc_hd__xor2_1 _07793_ (.A(_02041_),
    .B(_02042_),
    .X(_02089_));
 sky130_fd_sc_hd__a21o_1 _07794_ (.A1(_02088_),
    .A2(_02089_),
    .B1(_02043_),
    .X(_02090_));
 sky130_fd_sc_hd__xor2_1 _07795_ (.A(_02038_),
    .B(_02039_),
    .X(_02092_));
 sky130_fd_sc_hd__a21o_1 _07796_ (.A1(_02090_),
    .A2(_02092_),
    .B1(_02040_),
    .X(_02093_));
 sky130_fd_sc_hd__xor2_1 _07797_ (.A(_02034_),
    .B(_02035_),
    .X(_02094_));
 sky130_fd_sc_hd__a21oi_1 _07798_ (.A1(_02093_),
    .A2(_02094_),
    .B1(_02037_),
    .Y(_02095_));
 sky130_fd_sc_hd__nand2_1 _07799_ (.A(net36),
    .B(net25),
    .Y(_02096_));
 sky130_fd_sc_hd__and3_1 _07800_ (.A(_01963_),
    .B(_02026_),
    .C(_02096_),
    .X(_02097_));
 sky130_fd_sc_hd__and3_1 _07801_ (.A(net36),
    .B(net25),
    .C(_02027_),
    .X(_02098_));
 sky130_fd_sc_hd__o21ba_1 _07802_ (.A1(_02024_),
    .A2(_02033_),
    .B1_N(_02032_),
    .X(_02099_));
 sky130_fd_sc_hd__o21ai_1 _07803_ (.A1(_02097_),
    .A2(_02098_),
    .B1(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__nand2_1 _07804_ (.A(net37),
    .B(net24),
    .Y(_02101_));
 sky130_fd_sc_hd__and3_1 _07805_ (.A(net37),
    .B(net24),
    .C(_02100_),
    .X(_02103_));
 sky130_fd_sc_hd__xor2_1 _07806_ (.A(_02100_),
    .B(_02101_),
    .X(_02104_));
 sky130_fd_sc_hd__nor2_1 _07807_ (.A(_02095_),
    .B(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__xnor2_1 _07808_ (.A(_02095_),
    .B(_02104_),
    .Y(_02106_));
 sky130_fd_sc_hd__nand2_1 _07809_ (.A(net38),
    .B(net22),
    .Y(_02107_));
 sky130_fd_sc_hd__nor2_1 _07810_ (.A(_02106_),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__xnor2_1 _07811_ (.A(_02093_),
    .B(_02094_),
    .Y(_02109_));
 sky130_fd_sc_hd__nand2_1 _07812_ (.A(net38),
    .B(net21),
    .Y(_02110_));
 sky130_fd_sc_hd__nor2_1 _07813_ (.A(_02109_),
    .B(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__xnor2_1 _07814_ (.A(_02090_),
    .B(_02092_),
    .Y(_02112_));
 sky130_fd_sc_hd__nand2_1 _07815_ (.A(net38),
    .B(net20),
    .Y(_02114_));
 sky130_fd_sc_hd__nor2_1 _07816_ (.A(_02112_),
    .B(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__xnor2_1 _07817_ (.A(_02088_),
    .B(_02089_),
    .Y(_02116_));
 sky130_fd_sc_hd__nand2_1 _07818_ (.A(net38),
    .B(net19),
    .Y(_02117_));
 sky130_fd_sc_hd__nor2_1 _07819_ (.A(_02116_),
    .B(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__xnor2_1 _07820_ (.A(_02086_),
    .B(_02087_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_1 _07821_ (.A(net38),
    .B(net18),
    .Y(_02120_));
 sky130_fd_sc_hd__nor2_1 _07822_ (.A(_02119_),
    .B(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__xnor2_1 _07823_ (.A(_02084_),
    .B(_02085_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_1 _07824_ (.A(net38),
    .B(net17),
    .Y(_02123_));
 sky130_fd_sc_hd__nor2_1 _07825_ (.A(_02122_),
    .B(_02123_),
    .Y(_02125_));
 sky130_fd_sc_hd__xnor2_1 _07826_ (.A(_02082_),
    .B(_02083_),
    .Y(_02126_));
 sky130_fd_sc_hd__nand2_1 _07827_ (.A(net38),
    .B(net16),
    .Y(_02127_));
 sky130_fd_sc_hd__nor2_1 _07828_ (.A(_02126_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__xnor2_1 _07829_ (.A(_02079_),
    .B(_02081_),
    .Y(_02129_));
 sky130_fd_sc_hd__nand2_1 _07830_ (.A(net38),
    .B(net15),
    .Y(_02130_));
 sky130_fd_sc_hd__nor2_1 _07831_ (.A(_02129_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__xnor2_1 _07832_ (.A(_02077_),
    .B(_02078_),
    .Y(_02132_));
 sky130_fd_sc_hd__nand2_1 _07833_ (.A(net38),
    .B(net14),
    .Y(_02133_));
 sky130_fd_sc_hd__nor2_1 _07834_ (.A(_02132_),
    .B(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__xnor2_1 _07835_ (.A(_02075_),
    .B(_02076_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_1 _07836_ (.A(net38),
    .B(net13),
    .Y(_02137_));
 sky130_fd_sc_hd__nor2_1 _07837_ (.A(_02136_),
    .B(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__xnor2_1 _07838_ (.A(_02073_),
    .B(_02074_),
    .Y(_02139_));
 sky130_fd_sc_hd__nand2_1 _07839_ (.A(net38),
    .B(net11),
    .Y(_02140_));
 sky130_fd_sc_hd__nor2_1 _07840_ (.A(_02139_),
    .B(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__xnor2_1 _07841_ (.A(_02071_),
    .B(_02072_),
    .Y(_02142_));
 sky130_fd_sc_hd__nand2_1 _07842_ (.A(net38),
    .B(net10),
    .Y(_02143_));
 sky130_fd_sc_hd__nor2_1 _07843_ (.A(_02142_),
    .B(_02143_),
    .Y(_02144_));
 sky130_fd_sc_hd__a21o_1 _07844_ (.A1(_01503_),
    .A2(_01579_),
    .B1(_01578_),
    .X(_02145_));
 sky130_fd_sc_hd__xor2_1 _07845_ (.A(_02142_),
    .B(_02143_),
    .X(_02147_));
 sky130_fd_sc_hd__a21o_1 _07846_ (.A1(_02145_),
    .A2(_02147_),
    .B1(_02144_),
    .X(_02148_));
 sky130_fd_sc_hd__xor2_1 _07847_ (.A(_02139_),
    .B(_02140_),
    .X(_02149_));
 sky130_fd_sc_hd__a21o_1 _07848_ (.A1(_02148_),
    .A2(_02149_),
    .B1(_02141_),
    .X(_02150_));
 sky130_fd_sc_hd__xor2_1 _07849_ (.A(_02136_),
    .B(_02137_),
    .X(_02151_));
 sky130_fd_sc_hd__a21o_1 _07850_ (.A1(_02150_),
    .A2(_02151_),
    .B1(_02138_),
    .X(_02152_));
 sky130_fd_sc_hd__xor2_1 _07851_ (.A(_02132_),
    .B(_02133_),
    .X(_02153_));
 sky130_fd_sc_hd__a21o_1 _07852_ (.A1(_02152_),
    .A2(_02153_),
    .B1(_02134_),
    .X(_02154_));
 sky130_fd_sc_hd__xor2_1 _07853_ (.A(_02129_),
    .B(_02130_),
    .X(_02155_));
 sky130_fd_sc_hd__a21o_1 _07854_ (.A1(_02154_),
    .A2(_02155_),
    .B1(_02131_),
    .X(_02156_));
 sky130_fd_sc_hd__xor2_1 _07855_ (.A(_02126_),
    .B(_02127_),
    .X(_02158_));
 sky130_fd_sc_hd__a21o_1 _07856_ (.A1(_02156_),
    .A2(_02158_),
    .B1(_02128_),
    .X(_02159_));
 sky130_fd_sc_hd__xor2_1 _07857_ (.A(_02122_),
    .B(_02123_),
    .X(_02160_));
 sky130_fd_sc_hd__a21o_1 _07858_ (.A1(_02159_),
    .A2(_02160_),
    .B1(_02125_),
    .X(_02161_));
 sky130_fd_sc_hd__xor2_1 _07859_ (.A(_02119_),
    .B(_02120_),
    .X(_02162_));
 sky130_fd_sc_hd__a21o_1 _07860_ (.A1(_02161_),
    .A2(_02162_),
    .B1(_02121_),
    .X(_02163_));
 sky130_fd_sc_hd__xor2_1 _07861_ (.A(_02116_),
    .B(_02117_),
    .X(_02164_));
 sky130_fd_sc_hd__a21o_1 _07862_ (.A1(_02163_),
    .A2(_02164_),
    .B1(_02118_),
    .X(_02165_));
 sky130_fd_sc_hd__xor2_1 _07863_ (.A(_02112_),
    .B(_02114_),
    .X(_02166_));
 sky130_fd_sc_hd__a21o_1 _07864_ (.A1(_02165_),
    .A2(_02166_),
    .B1(_02115_),
    .X(_02167_));
 sky130_fd_sc_hd__xor2_1 _07865_ (.A(_02109_),
    .B(_02110_),
    .X(_02169_));
 sky130_fd_sc_hd__a21o_1 _07866_ (.A1(_02167_),
    .A2(_02169_),
    .B1(_02111_),
    .X(_02170_));
 sky130_fd_sc_hd__xor2_1 _07867_ (.A(_02106_),
    .B(_02107_),
    .X(_02171_));
 sky130_fd_sc_hd__a21oi_1 _07868_ (.A1(_02170_),
    .A2(_02171_),
    .B1(_02108_),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _07869_ (.A(net37),
    .B(net25),
    .Y(_02173_));
 sky130_fd_sc_hd__nand2_1 _07870_ (.A(_02097_),
    .B(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__or2_1 _07871_ (.A(_02097_),
    .B(_02173_),
    .X(_02175_));
 sky130_fd_sc_hd__a211o_1 _07872_ (.A1(_02174_),
    .A2(_02175_),
    .B1(_02103_),
    .C1(_02105_),
    .X(_02176_));
 sky130_fd_sc_hd__nand2_1 _07873_ (.A(net38),
    .B(net24),
    .Y(_02177_));
 sky130_fd_sc_hd__and3_1 _07874_ (.A(net38),
    .B(net24),
    .C(_02176_),
    .X(_02178_));
 sky130_fd_sc_hd__xor2_1 _07875_ (.A(_02176_),
    .B(_02177_),
    .X(_02180_));
 sky130_fd_sc_hd__xnor2_1 _07876_ (.A(_02172_),
    .B(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _07877_ (.A(net39),
    .B(net22),
    .Y(_02182_));
 sky130_fd_sc_hd__nor2_1 _07878_ (.A(_02181_),
    .B(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__xnor2_1 _07879_ (.A(_02170_),
    .B(_02171_),
    .Y(_02184_));
 sky130_fd_sc_hd__nand2_1 _07880_ (.A(net39),
    .B(net21),
    .Y(_02185_));
 sky130_fd_sc_hd__nor2_1 _07881_ (.A(_02184_),
    .B(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__xnor2_1 _07882_ (.A(_02167_),
    .B(_02169_),
    .Y(_02187_));
 sky130_fd_sc_hd__nand2_1 _07883_ (.A(net39),
    .B(net20),
    .Y(_02188_));
 sky130_fd_sc_hd__nor2_1 _07884_ (.A(_02187_),
    .B(_02188_),
    .Y(_02189_));
 sky130_fd_sc_hd__xnor2_1 _07885_ (.A(_02165_),
    .B(_02166_),
    .Y(_02191_));
 sky130_fd_sc_hd__nand2_1 _07886_ (.A(net39),
    .B(net19),
    .Y(_02192_));
 sky130_fd_sc_hd__nor2_1 _07887_ (.A(_02191_),
    .B(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__xnor2_1 _07888_ (.A(_02163_),
    .B(_02164_),
    .Y(_02194_));
 sky130_fd_sc_hd__nand2_1 _07889_ (.A(net39),
    .B(net18),
    .Y(_02195_));
 sky130_fd_sc_hd__nor2_1 _07890_ (.A(_02194_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__xnor2_1 _07891_ (.A(_02161_),
    .B(_02162_),
    .Y(_02197_));
 sky130_fd_sc_hd__nand2_1 _07892_ (.A(net39),
    .B(net17),
    .Y(_02198_));
 sky130_fd_sc_hd__nor2_1 _07893_ (.A(_02197_),
    .B(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__xnor2_1 _07894_ (.A(_02159_),
    .B(_02160_),
    .Y(_02200_));
 sky130_fd_sc_hd__nand2_1 _07895_ (.A(net39),
    .B(net16),
    .Y(_02202_));
 sky130_fd_sc_hd__nor2_1 _07896_ (.A(_02200_),
    .B(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__xnor2_1 _07897_ (.A(_02156_),
    .B(_02158_),
    .Y(_02204_));
 sky130_fd_sc_hd__nand2_1 _07898_ (.A(net39),
    .B(net15),
    .Y(_02205_));
 sky130_fd_sc_hd__nor2_1 _07899_ (.A(_02204_),
    .B(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__xnor2_1 _07900_ (.A(_02154_),
    .B(_02155_),
    .Y(_02207_));
 sky130_fd_sc_hd__nand2_1 _07901_ (.A(net39),
    .B(net14),
    .Y(_02208_));
 sky130_fd_sc_hd__nor2_1 _07902_ (.A(_02207_),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__xnor2_1 _07903_ (.A(_02152_),
    .B(_02153_),
    .Y(_02210_));
 sky130_fd_sc_hd__nand2_1 _07904_ (.A(net39),
    .B(net13),
    .Y(_02211_));
 sky130_fd_sc_hd__nor2_1 _07905_ (.A(_02210_),
    .B(_02211_),
    .Y(_02213_));
 sky130_fd_sc_hd__xnor2_1 _07906_ (.A(_02150_),
    .B(_02151_),
    .Y(_02214_));
 sky130_fd_sc_hd__nand2_1 _07907_ (.A(net39),
    .B(net11),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _07908_ (.A(_02214_),
    .B(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__xnor2_1 _07909_ (.A(_02148_),
    .B(_02149_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_1 _07910_ (.A(net39),
    .B(net10),
    .Y(_02218_));
 sky130_fd_sc_hd__nor2_1 _07911_ (.A(_02217_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__xnor2_1 _07912_ (.A(_02145_),
    .B(_02147_),
    .Y(_02220_));
 sky130_fd_sc_hd__nand2_1 _07913_ (.A(net39),
    .B(net9),
    .Y(_02221_));
 sky130_fd_sc_hd__nor2_1 _07914_ (.A(_02220_),
    .B(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__a21o_1 _07915_ (.A1(_01501_),
    .A2(_01582_),
    .B1(_01581_),
    .X(_02224_));
 sky130_fd_sc_hd__xor2_1 _07916_ (.A(_02220_),
    .B(_02221_),
    .X(_02225_));
 sky130_fd_sc_hd__a21o_1 _07917_ (.A1(_02224_),
    .A2(_02225_),
    .B1(_02222_),
    .X(_02226_));
 sky130_fd_sc_hd__xor2_1 _07918_ (.A(_02217_),
    .B(_02218_),
    .X(_02227_));
 sky130_fd_sc_hd__a21o_1 _07919_ (.A1(_02226_),
    .A2(_02227_),
    .B1(_02219_),
    .X(_02228_));
 sky130_fd_sc_hd__xor2_1 _07920_ (.A(_02214_),
    .B(_02215_),
    .X(_02229_));
 sky130_fd_sc_hd__a21o_1 _07921_ (.A1(_02228_),
    .A2(_02229_),
    .B1(_02216_),
    .X(_02230_));
 sky130_fd_sc_hd__xor2_1 _07922_ (.A(_02210_),
    .B(_02211_),
    .X(_02231_));
 sky130_fd_sc_hd__a21o_1 _07923_ (.A1(_02230_),
    .A2(_02231_),
    .B1(_02213_),
    .X(_02232_));
 sky130_fd_sc_hd__xor2_1 _07924_ (.A(_02207_),
    .B(_02208_),
    .X(_02233_));
 sky130_fd_sc_hd__a21o_1 _07925_ (.A1(_02232_),
    .A2(_02233_),
    .B1(_02209_),
    .X(_02235_));
 sky130_fd_sc_hd__xor2_1 _07926_ (.A(_02204_),
    .B(_02205_),
    .X(_02236_));
 sky130_fd_sc_hd__a21o_1 _07927_ (.A1(_02235_),
    .A2(_02236_),
    .B1(_02206_),
    .X(_02237_));
 sky130_fd_sc_hd__xor2_1 _07928_ (.A(_02200_),
    .B(_02202_),
    .X(_02238_));
 sky130_fd_sc_hd__a21o_1 _07929_ (.A1(_02237_),
    .A2(_02238_),
    .B1(_02203_),
    .X(_02239_));
 sky130_fd_sc_hd__xor2_1 _07930_ (.A(_02197_),
    .B(_02198_),
    .X(_02240_));
 sky130_fd_sc_hd__a21o_1 _07931_ (.A1(_02239_),
    .A2(_02240_),
    .B1(_02199_),
    .X(_02241_));
 sky130_fd_sc_hd__xor2_1 _07932_ (.A(_02194_),
    .B(_02195_),
    .X(_02242_));
 sky130_fd_sc_hd__a21o_1 _07933_ (.A1(_02241_),
    .A2(_02242_),
    .B1(_02196_),
    .X(_02243_));
 sky130_fd_sc_hd__xor2_1 _07934_ (.A(_02191_),
    .B(_02192_),
    .X(_02244_));
 sky130_fd_sc_hd__a21o_1 _07935_ (.A1(_02243_),
    .A2(_02244_),
    .B1(_02193_),
    .X(_02246_));
 sky130_fd_sc_hd__xor2_1 _07936_ (.A(_02187_),
    .B(_02188_),
    .X(_02247_));
 sky130_fd_sc_hd__a21o_1 _07937_ (.A1(_02246_),
    .A2(_02247_),
    .B1(_02189_),
    .X(_02248_));
 sky130_fd_sc_hd__xor2_1 _07938_ (.A(_02184_),
    .B(_02185_),
    .X(_02249_));
 sky130_fd_sc_hd__a21o_1 _07939_ (.A1(_02248_),
    .A2(_02249_),
    .B1(_02186_),
    .X(_02250_));
 sky130_fd_sc_hd__xor2_1 _07940_ (.A(_02181_),
    .B(_02182_),
    .X(_02251_));
 sky130_fd_sc_hd__a21oi_1 _07941_ (.A1(_02250_),
    .A2(_02251_),
    .B1(_02183_),
    .Y(_02252_));
 sky130_fd_sc_hd__nand2_1 _07942_ (.A(net38),
    .B(net25),
    .Y(_02253_));
 sky130_fd_sc_hd__and3_1 _07943_ (.A(_02097_),
    .B(_02173_),
    .C(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__and3_1 _07944_ (.A(net38),
    .B(net25),
    .C(_02174_),
    .X(_02255_));
 sky130_fd_sc_hd__o21ba_1 _07945_ (.A1(_02172_),
    .A2(_02180_),
    .B1_N(_02178_),
    .X(_02257_));
 sky130_fd_sc_hd__o21ai_1 _07946_ (.A1(_02254_),
    .A2(_02255_),
    .B1(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__nand2_1 _07947_ (.A(net39),
    .B(net24),
    .Y(_02259_));
 sky130_fd_sc_hd__xor2_1 _07948_ (.A(_02258_),
    .B(_02259_),
    .X(_02260_));
 sky130_fd_sc_hd__xnor2_1 _07949_ (.A(_02252_),
    .B(_02260_),
    .Y(_02261_));
 sky130_fd_sc_hd__nand2_1 _07950_ (.A(net40),
    .B(net22),
    .Y(_02262_));
 sky130_fd_sc_hd__nor2_1 _07951_ (.A(_02261_),
    .B(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__xnor2_1 _07952_ (.A(_02250_),
    .B(_02251_),
    .Y(_02264_));
 sky130_fd_sc_hd__nand2_1 _07953_ (.A(net40),
    .B(net21),
    .Y(_02265_));
 sky130_fd_sc_hd__nor2_1 _07954_ (.A(_02264_),
    .B(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__xnor2_1 _07955_ (.A(_02248_),
    .B(_02249_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand2_1 _07956_ (.A(net40),
    .B(net20),
    .Y(_02269_));
 sky130_fd_sc_hd__nor2_1 _07957_ (.A(_02268_),
    .B(_02269_),
    .Y(_02270_));
 sky130_fd_sc_hd__xnor2_1 _07958_ (.A(_02246_),
    .B(_02247_),
    .Y(_02271_));
 sky130_fd_sc_hd__nand2_1 _07959_ (.A(net40),
    .B(net19),
    .Y(_02272_));
 sky130_fd_sc_hd__nor2_1 _07960_ (.A(_02271_),
    .B(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hd__xnor2_1 _07961_ (.A(_02243_),
    .B(_02244_),
    .Y(_02274_));
 sky130_fd_sc_hd__nand2_1 _07962_ (.A(net40),
    .B(net18),
    .Y(_02275_));
 sky130_fd_sc_hd__nor2_1 _07963_ (.A(_02274_),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__xnor2_1 _07964_ (.A(_02241_),
    .B(_02242_),
    .Y(_02277_));
 sky130_fd_sc_hd__nand2_1 _07965_ (.A(net40),
    .B(net17),
    .Y(_02279_));
 sky130_fd_sc_hd__nor2_1 _07966_ (.A(_02277_),
    .B(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__xnor2_1 _07967_ (.A(_02239_),
    .B(_02240_),
    .Y(_02281_));
 sky130_fd_sc_hd__nand2_1 _07968_ (.A(net40),
    .B(net16),
    .Y(_02282_));
 sky130_fd_sc_hd__nor2_1 _07969_ (.A(_02281_),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__xnor2_1 _07970_ (.A(_02237_),
    .B(_02238_),
    .Y(_02284_));
 sky130_fd_sc_hd__nand2_1 _07971_ (.A(net40),
    .B(net15),
    .Y(_02285_));
 sky130_fd_sc_hd__nor2_1 _07972_ (.A(_02284_),
    .B(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hd__xnor2_1 _07973_ (.A(_02235_),
    .B(_02236_),
    .Y(_02287_));
 sky130_fd_sc_hd__nand2_1 _07974_ (.A(net40),
    .B(net14),
    .Y(_02288_));
 sky130_fd_sc_hd__nor2_1 _07975_ (.A(_02287_),
    .B(_02288_),
    .Y(_02290_));
 sky130_fd_sc_hd__xnor2_1 _07976_ (.A(_02232_),
    .B(_02233_),
    .Y(_02291_));
 sky130_fd_sc_hd__nand2_1 _07977_ (.A(net40),
    .B(net13),
    .Y(_02292_));
 sky130_fd_sc_hd__nor2_1 _07978_ (.A(_02291_),
    .B(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__xnor2_1 _07979_ (.A(_02230_),
    .B(_02231_),
    .Y(_02294_));
 sky130_fd_sc_hd__nand2_1 _07980_ (.A(net40),
    .B(net11),
    .Y(_02295_));
 sky130_fd_sc_hd__nor2_1 _07981_ (.A(_02294_),
    .B(_02295_),
    .Y(_02296_));
 sky130_fd_sc_hd__xnor2_1 _07982_ (.A(_02228_),
    .B(_02229_),
    .Y(_02297_));
 sky130_fd_sc_hd__nand2_1 _07983_ (.A(net40),
    .B(net10),
    .Y(_02298_));
 sky130_fd_sc_hd__nor2_1 _07984_ (.A(_02297_),
    .B(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__xnor2_1 _07985_ (.A(_02226_),
    .B(_02227_),
    .Y(_02301_));
 sky130_fd_sc_hd__nand2_1 _07986_ (.A(net40),
    .B(net9),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_1 _07987_ (.A(_02301_),
    .B(_02302_),
    .Y(_02303_));
 sky130_fd_sc_hd__xnor2_1 _07988_ (.A(_02224_),
    .B(_02225_),
    .Y(_02304_));
 sky130_fd_sc_hd__nand2_1 _07989_ (.A(net8),
    .B(net40),
    .Y(_02305_));
 sky130_fd_sc_hd__nor2_1 _07990_ (.A(_02304_),
    .B(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__a21o_1 _07991_ (.A1(_01499_),
    .A2(_01585_),
    .B1(_01584_),
    .X(_02307_));
 sky130_fd_sc_hd__xor2_1 _07992_ (.A(_02304_),
    .B(_02305_),
    .X(_02308_));
 sky130_fd_sc_hd__a21o_1 _07993_ (.A1(_02307_),
    .A2(_02308_),
    .B1(_02306_),
    .X(_02309_));
 sky130_fd_sc_hd__xor2_1 _07994_ (.A(_02301_),
    .B(_02302_),
    .X(_02310_));
 sky130_fd_sc_hd__a21o_1 _07995_ (.A1(_02309_),
    .A2(_02310_),
    .B1(_02303_),
    .X(_02312_));
 sky130_fd_sc_hd__xor2_1 _07996_ (.A(_02297_),
    .B(_02298_),
    .X(_02313_));
 sky130_fd_sc_hd__a21o_1 _07997_ (.A1(_02312_),
    .A2(_02313_),
    .B1(_02299_),
    .X(_02314_));
 sky130_fd_sc_hd__xor2_1 _07998_ (.A(_02294_),
    .B(_02295_),
    .X(_02315_));
 sky130_fd_sc_hd__a21o_1 _07999_ (.A1(_02314_),
    .A2(_02315_),
    .B1(_02296_),
    .X(_02316_));
 sky130_fd_sc_hd__xor2_1 _08000_ (.A(_02291_),
    .B(_02292_),
    .X(_02317_));
 sky130_fd_sc_hd__a21o_1 _08001_ (.A1(_02316_),
    .A2(_02317_),
    .B1(_02293_),
    .X(_02318_));
 sky130_fd_sc_hd__xor2_1 _08002_ (.A(_02287_),
    .B(_02288_),
    .X(_02319_));
 sky130_fd_sc_hd__a21o_1 _08003_ (.A1(_02318_),
    .A2(_02319_),
    .B1(_02290_),
    .X(_02320_));
 sky130_fd_sc_hd__xor2_1 _08004_ (.A(_02284_),
    .B(_02285_),
    .X(_02321_));
 sky130_fd_sc_hd__a21o_1 _08005_ (.A1(_02320_),
    .A2(_02321_),
    .B1(_02286_),
    .X(_02323_));
 sky130_fd_sc_hd__xor2_1 _08006_ (.A(_02281_),
    .B(_02282_),
    .X(_02324_));
 sky130_fd_sc_hd__a21o_1 _08007_ (.A1(_02323_),
    .A2(_02324_),
    .B1(_02283_),
    .X(_02325_));
 sky130_fd_sc_hd__xor2_1 _08008_ (.A(_02277_),
    .B(_02279_),
    .X(_02326_));
 sky130_fd_sc_hd__a21o_1 _08009_ (.A1(_02325_),
    .A2(_02326_),
    .B1(_02280_),
    .X(_02327_));
 sky130_fd_sc_hd__xor2_1 _08010_ (.A(_02274_),
    .B(_02275_),
    .X(_02328_));
 sky130_fd_sc_hd__a21o_1 _08011_ (.A1(_02327_),
    .A2(_02328_),
    .B1(_02276_),
    .X(_02329_));
 sky130_fd_sc_hd__xor2_1 _08012_ (.A(_02271_),
    .B(_02272_),
    .X(_02330_));
 sky130_fd_sc_hd__a21o_1 _08013_ (.A1(_02329_),
    .A2(_02330_),
    .B1(_02273_),
    .X(_02331_));
 sky130_fd_sc_hd__xor2_1 _08014_ (.A(_02268_),
    .B(_02269_),
    .X(_02332_));
 sky130_fd_sc_hd__a21o_1 _08015_ (.A1(_02331_),
    .A2(_02332_),
    .B1(_02270_),
    .X(_02334_));
 sky130_fd_sc_hd__xor2_1 _08016_ (.A(_02264_),
    .B(_02265_),
    .X(_02335_));
 sky130_fd_sc_hd__a21o_1 _08017_ (.A1(_02334_),
    .A2(_02335_),
    .B1(_02266_),
    .X(_02336_));
 sky130_fd_sc_hd__xor2_1 _08018_ (.A(_02261_),
    .B(_02262_),
    .X(_02337_));
 sky130_fd_sc_hd__a21oi_1 _08019_ (.A1(_02336_),
    .A2(_02337_),
    .B1(_02263_),
    .Y(_02338_));
 sky130_fd_sc_hd__nand2_1 _08020_ (.A(net39),
    .B(net25),
    .Y(_02339_));
 sky130_fd_sc_hd__and2_1 _08021_ (.A(_02254_),
    .B(_02339_),
    .X(_02340_));
 sky130_fd_sc_hd__nor2_1 _08022_ (.A(_02254_),
    .B(_02339_),
    .Y(_02341_));
 sky130_fd_sc_hd__o22ai_1 _08023_ (.A1(_02252_),
    .A2(_02260_),
    .B1(_02340_),
    .B2(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hd__a31o_1 _08024_ (.A1(net39),
    .A2(net24),
    .A3(_02258_),
    .B1(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__nand2_1 _08025_ (.A(net40),
    .B(net24),
    .Y(_02345_));
 sky130_fd_sc_hd__xor2_1 _08026_ (.A(_02343_),
    .B(_02345_),
    .X(_02346_));
 sky130_fd_sc_hd__xnor2_1 _08027_ (.A(_02338_),
    .B(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_1 _08028_ (.A(net41),
    .B(net22),
    .Y(_02348_));
 sky130_fd_sc_hd__nor2_1 _08029_ (.A(_02347_),
    .B(_02348_),
    .Y(_02349_));
 sky130_fd_sc_hd__xnor2_1 _08030_ (.A(_02336_),
    .B(_02337_),
    .Y(_02350_));
 sky130_fd_sc_hd__nand2_1 _08031_ (.A(net41),
    .B(net21),
    .Y(_02351_));
 sky130_fd_sc_hd__nor2_1 _08032_ (.A(_02350_),
    .B(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__xnor2_1 _08033_ (.A(_02334_),
    .B(_02335_),
    .Y(_02353_));
 sky130_fd_sc_hd__nand2_1 _08034_ (.A(net41),
    .B(net20),
    .Y(_02354_));
 sky130_fd_sc_hd__nor2_1 _08035_ (.A(_02353_),
    .B(_02354_),
    .Y(_02356_));
 sky130_fd_sc_hd__xnor2_1 _08036_ (.A(_02331_),
    .B(_02332_),
    .Y(_02357_));
 sky130_fd_sc_hd__nand2_1 _08037_ (.A(net41),
    .B(net19),
    .Y(_02358_));
 sky130_fd_sc_hd__nor2_1 _08038_ (.A(_02357_),
    .B(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__xnor2_1 _08039_ (.A(_02329_),
    .B(_02330_),
    .Y(_02360_));
 sky130_fd_sc_hd__nand2_1 _08040_ (.A(net41),
    .B(net18),
    .Y(_02361_));
 sky130_fd_sc_hd__nor2_1 _08041_ (.A(_02360_),
    .B(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__xnor2_1 _08042_ (.A(_02327_),
    .B(_02328_),
    .Y(_02363_));
 sky130_fd_sc_hd__nand2_1 _08043_ (.A(net41),
    .B(net17),
    .Y(_02364_));
 sky130_fd_sc_hd__nor2_1 _08044_ (.A(_02363_),
    .B(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__xnor2_1 _08045_ (.A(_02325_),
    .B(_02326_),
    .Y(_02367_));
 sky130_fd_sc_hd__nand2_1 _08046_ (.A(net41),
    .B(net16),
    .Y(_02368_));
 sky130_fd_sc_hd__nor2_1 _08047_ (.A(_02367_),
    .B(_02368_),
    .Y(_02369_));
 sky130_fd_sc_hd__xnor2_1 _08048_ (.A(_02323_),
    .B(_02324_),
    .Y(_02370_));
 sky130_fd_sc_hd__nand2_1 _08049_ (.A(net41),
    .B(net15),
    .Y(_02371_));
 sky130_fd_sc_hd__nor2_1 _08050_ (.A(_02370_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__xnor2_1 _08051_ (.A(_02320_),
    .B(_02321_),
    .Y(_02373_));
 sky130_fd_sc_hd__nand2_1 _08052_ (.A(net41),
    .B(net14),
    .Y(_02374_));
 sky130_fd_sc_hd__nor2_1 _08053_ (.A(_02373_),
    .B(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__xnor2_1 _08054_ (.A(_02318_),
    .B(_02319_),
    .Y(_02376_));
 sky130_fd_sc_hd__nand2_1 _08055_ (.A(net41),
    .B(net13),
    .Y(_02378_));
 sky130_fd_sc_hd__nor2_1 _08056_ (.A(_02376_),
    .B(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__xnor2_1 _08057_ (.A(_02316_),
    .B(_02317_),
    .Y(_02380_));
 sky130_fd_sc_hd__nand2_1 _08058_ (.A(net41),
    .B(net11),
    .Y(_02381_));
 sky130_fd_sc_hd__nor2_1 _08059_ (.A(_02380_),
    .B(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__xnor2_1 _08060_ (.A(_02314_),
    .B(_02315_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand2_1 _08061_ (.A(net41),
    .B(net10),
    .Y(_02384_));
 sky130_fd_sc_hd__nor2_1 _08062_ (.A(_02383_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__xnor2_1 _08063_ (.A(_02312_),
    .B(_02313_),
    .Y(_02386_));
 sky130_fd_sc_hd__nand2_1 _08064_ (.A(net9),
    .B(net41),
    .Y(_02387_));
 sky130_fd_sc_hd__nor2_1 _08065_ (.A(_02386_),
    .B(_02387_),
    .Y(_02389_));
 sky130_fd_sc_hd__xnor2_1 _08066_ (.A(_02309_),
    .B(_02310_),
    .Y(_02390_));
 sky130_fd_sc_hd__nand2_1 _08067_ (.A(net8),
    .B(net41),
    .Y(_02391_));
 sky130_fd_sc_hd__nor2_1 _08068_ (.A(_02390_),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__xnor2_1 _08069_ (.A(_02307_),
    .B(_02308_),
    .Y(_02393_));
 sky130_fd_sc_hd__nand2_1 _08070_ (.A(net7),
    .B(net41),
    .Y(_02394_));
 sky130_fd_sc_hd__nor2_1 _08071_ (.A(_02393_),
    .B(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__a21o_1 _08072_ (.A1(_01496_),
    .A2(_01589_),
    .B1(_01588_),
    .X(_02396_));
 sky130_fd_sc_hd__xor2_1 _08073_ (.A(_02393_),
    .B(_02394_),
    .X(_02397_));
 sky130_fd_sc_hd__a21o_1 _08074_ (.A1(_02396_),
    .A2(_02397_),
    .B1(_02395_),
    .X(_02398_));
 sky130_fd_sc_hd__xor2_1 _08075_ (.A(_02390_),
    .B(_02391_),
    .X(_02400_));
 sky130_fd_sc_hd__a21o_1 _08076_ (.A1(_02398_),
    .A2(_02400_),
    .B1(_02392_),
    .X(_02401_));
 sky130_fd_sc_hd__xor2_1 _08077_ (.A(_02386_),
    .B(_02387_),
    .X(_02402_));
 sky130_fd_sc_hd__a21o_1 _08078_ (.A1(_02401_),
    .A2(_02402_),
    .B1(_02389_),
    .X(_02403_));
 sky130_fd_sc_hd__xor2_1 _08079_ (.A(_02383_),
    .B(_02384_),
    .X(_02404_));
 sky130_fd_sc_hd__a21o_1 _08080_ (.A1(_02403_),
    .A2(_02404_),
    .B1(_02385_),
    .X(_02405_));
 sky130_fd_sc_hd__xor2_1 _08081_ (.A(_02380_),
    .B(_02381_),
    .X(_02406_));
 sky130_fd_sc_hd__a21o_1 _08082_ (.A1(_02405_),
    .A2(_02406_),
    .B1(_02382_),
    .X(_02407_));
 sky130_fd_sc_hd__xor2_1 _08083_ (.A(_02376_),
    .B(_02378_),
    .X(_02408_));
 sky130_fd_sc_hd__a21o_1 _08084_ (.A1(_02407_),
    .A2(_02408_),
    .B1(_02379_),
    .X(_02409_));
 sky130_fd_sc_hd__xor2_1 _08085_ (.A(_02373_),
    .B(_02374_),
    .X(_02411_));
 sky130_fd_sc_hd__a21o_1 _08086_ (.A1(_02409_),
    .A2(_02411_),
    .B1(_02375_),
    .X(_02412_));
 sky130_fd_sc_hd__xor2_1 _08087_ (.A(_02370_),
    .B(_02371_),
    .X(_02413_));
 sky130_fd_sc_hd__a21o_1 _08088_ (.A1(_02412_),
    .A2(_02413_),
    .B1(_02372_),
    .X(_02414_));
 sky130_fd_sc_hd__xor2_1 _08089_ (.A(_02367_),
    .B(_02368_),
    .X(_02415_));
 sky130_fd_sc_hd__a21o_1 _08090_ (.A1(_02414_),
    .A2(_02415_),
    .B1(_02369_),
    .X(_02416_));
 sky130_fd_sc_hd__xor2_1 _08091_ (.A(_02363_),
    .B(_02364_),
    .X(_02417_));
 sky130_fd_sc_hd__a21o_1 _08092_ (.A1(_02416_),
    .A2(_02417_),
    .B1(_02365_),
    .X(_02418_));
 sky130_fd_sc_hd__xor2_1 _08093_ (.A(_02360_),
    .B(_02361_),
    .X(_02419_));
 sky130_fd_sc_hd__a21o_1 _08094_ (.A1(_02418_),
    .A2(_02419_),
    .B1(_02362_),
    .X(_02420_));
 sky130_fd_sc_hd__xor2_1 _08095_ (.A(_02357_),
    .B(_02358_),
    .X(_02422_));
 sky130_fd_sc_hd__a21o_1 _08096_ (.A1(_02420_),
    .A2(_02422_),
    .B1(_02359_),
    .X(_02423_));
 sky130_fd_sc_hd__xor2_1 _08097_ (.A(_02353_),
    .B(_02354_),
    .X(_02424_));
 sky130_fd_sc_hd__a21o_1 _08098_ (.A1(_02423_),
    .A2(_02424_),
    .B1(_02356_),
    .X(_02425_));
 sky130_fd_sc_hd__xor2_1 _08099_ (.A(_02350_),
    .B(_02351_),
    .X(_02426_));
 sky130_fd_sc_hd__a21o_1 _08100_ (.A1(_02425_),
    .A2(_02426_),
    .B1(_02352_),
    .X(_02427_));
 sky130_fd_sc_hd__xor2_1 _08101_ (.A(_02347_),
    .B(_02348_),
    .X(_02428_));
 sky130_fd_sc_hd__a21oi_1 _08102_ (.A1(_02427_),
    .A2(_02428_),
    .B1(_02349_),
    .Y(_02429_));
 sky130_fd_sc_hd__nand2_1 _08103_ (.A(net40),
    .B(net25),
    .Y(_02430_));
 sky130_fd_sc_hd__nand2_1 _08104_ (.A(_02340_),
    .B(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__or2_1 _08105_ (.A(_02340_),
    .B(_02430_),
    .X(_02433_));
 sky130_fd_sc_hd__a2bb2o_1 _08106_ (.A1_N(_02338_),
    .A2_N(_02346_),
    .B1(_02431_),
    .B2(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__a31o_1 _08107_ (.A1(net40),
    .A2(net24),
    .A3(_02343_),
    .B1(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__nand2_1 _08108_ (.A(net41),
    .B(net24),
    .Y(_02436_));
 sky130_fd_sc_hd__xor2_1 _08109_ (.A(_02435_),
    .B(_02436_),
    .X(_02437_));
 sky130_fd_sc_hd__nor2_1 _08110_ (.A(_02429_),
    .B(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__xnor2_1 _08111_ (.A(_02429_),
    .B(_02437_),
    .Y(_02439_));
 sky130_fd_sc_hd__nand2_1 _08112_ (.A(net42),
    .B(net22),
    .Y(_02440_));
 sky130_fd_sc_hd__nor2_1 _08113_ (.A(_02439_),
    .B(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__xnor2_1 _08114_ (.A(_02427_),
    .B(_02428_),
    .Y(_02442_));
 sky130_fd_sc_hd__nand2_1 _08115_ (.A(net42),
    .B(net21),
    .Y(_02444_));
 sky130_fd_sc_hd__nor2_1 _08116_ (.A(_02442_),
    .B(_02444_),
    .Y(_02445_));
 sky130_fd_sc_hd__xnor2_1 _08117_ (.A(_02425_),
    .B(_02426_),
    .Y(_02446_));
 sky130_fd_sc_hd__nand2_1 _08118_ (.A(net42),
    .B(net20),
    .Y(_02447_));
 sky130_fd_sc_hd__nor2_1 _08119_ (.A(_02446_),
    .B(_02447_),
    .Y(_02448_));
 sky130_fd_sc_hd__xnor2_1 _08120_ (.A(_02423_),
    .B(_02424_),
    .Y(_02449_));
 sky130_fd_sc_hd__nand2_1 _08121_ (.A(net42),
    .B(net19),
    .Y(_02450_));
 sky130_fd_sc_hd__nor2_1 _08122_ (.A(_02449_),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__xnor2_1 _08123_ (.A(_02420_),
    .B(_02422_),
    .Y(_02452_));
 sky130_fd_sc_hd__nand2_1 _08124_ (.A(net42),
    .B(net18),
    .Y(_02453_));
 sky130_fd_sc_hd__nor2_1 _08125_ (.A(_02452_),
    .B(_02453_),
    .Y(_02455_));
 sky130_fd_sc_hd__xnor2_1 _08126_ (.A(_02418_),
    .B(_02419_),
    .Y(_02456_));
 sky130_fd_sc_hd__nand2_1 _08127_ (.A(net42),
    .B(net17),
    .Y(_02457_));
 sky130_fd_sc_hd__nor2_1 _08128_ (.A(_02456_),
    .B(_02457_),
    .Y(_02458_));
 sky130_fd_sc_hd__xnor2_1 _08129_ (.A(_02416_),
    .B(_02417_),
    .Y(_02459_));
 sky130_fd_sc_hd__nand2_1 _08130_ (.A(net42),
    .B(net16),
    .Y(_02460_));
 sky130_fd_sc_hd__nor2_1 _08131_ (.A(_02459_),
    .B(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__xnor2_1 _08132_ (.A(_02414_),
    .B(_02415_),
    .Y(_02462_));
 sky130_fd_sc_hd__nand2_1 _08133_ (.A(net42),
    .B(net15),
    .Y(_02463_));
 sky130_fd_sc_hd__nor2_1 _08134_ (.A(_02462_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__xnor2_1 _08135_ (.A(_02412_),
    .B(_02413_),
    .Y(_02466_));
 sky130_fd_sc_hd__nand2_1 _08136_ (.A(net42),
    .B(net14),
    .Y(_02467_));
 sky130_fd_sc_hd__nor2_1 _08137_ (.A(_02466_),
    .B(_02467_),
    .Y(_02468_));
 sky130_fd_sc_hd__xnor2_1 _08138_ (.A(_02409_),
    .B(_02411_),
    .Y(_02469_));
 sky130_fd_sc_hd__nand2_1 _08139_ (.A(net42),
    .B(net13),
    .Y(_02470_));
 sky130_fd_sc_hd__nor2_1 _08140_ (.A(_02469_),
    .B(_02470_),
    .Y(_02471_));
 sky130_fd_sc_hd__xnor2_1 _08141_ (.A(_02407_),
    .B(_02408_),
    .Y(_02472_));
 sky130_fd_sc_hd__nand2_1 _08142_ (.A(net42),
    .B(net11),
    .Y(_02473_));
 sky130_fd_sc_hd__nor2_1 _08143_ (.A(_02472_),
    .B(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__xnor2_1 _08144_ (.A(_02405_),
    .B(_02406_),
    .Y(_02475_));
 sky130_fd_sc_hd__nand2_1 _08145_ (.A(net10),
    .B(net42),
    .Y(_02477_));
 sky130_fd_sc_hd__nor2_1 _08146_ (.A(_02475_),
    .B(_02477_),
    .Y(_02478_));
 sky130_fd_sc_hd__xnor2_1 _08147_ (.A(_02403_),
    .B(_02404_),
    .Y(_02479_));
 sky130_fd_sc_hd__nand2_1 _08148_ (.A(net9),
    .B(net42),
    .Y(_02480_));
 sky130_fd_sc_hd__nor2_1 _08149_ (.A(_02479_),
    .B(_02480_),
    .Y(_02481_));
 sky130_fd_sc_hd__xnor2_1 _08150_ (.A(_02401_),
    .B(_02402_),
    .Y(_02482_));
 sky130_fd_sc_hd__nand2_1 _08151_ (.A(net8),
    .B(net42),
    .Y(_02483_));
 sky130_fd_sc_hd__nor2_1 _08152_ (.A(_02482_),
    .B(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__xnor2_1 _08153_ (.A(_02398_),
    .B(_02400_),
    .Y(_02485_));
 sky130_fd_sc_hd__nand2_1 _08154_ (.A(net7),
    .B(net42),
    .Y(_02486_));
 sky130_fd_sc_hd__nor2_1 _08155_ (.A(_02485_),
    .B(_02486_),
    .Y(_02488_));
 sky130_fd_sc_hd__xnor2_1 _08156_ (.A(_02396_),
    .B(_02397_),
    .Y(_02489_));
 sky130_fd_sc_hd__nand2_1 _08157_ (.A(net6),
    .B(net42),
    .Y(_02490_));
 sky130_fd_sc_hd__nor2_1 _08158_ (.A(_02489_),
    .B(_02490_),
    .Y(_02491_));
 sky130_fd_sc_hd__a21o_1 _08159_ (.A1(_01494_),
    .A2(_01592_),
    .B1(_01591_),
    .X(_02492_));
 sky130_fd_sc_hd__xor2_1 _08160_ (.A(_02489_),
    .B(_02490_),
    .X(_02493_));
 sky130_fd_sc_hd__a21o_1 _08161_ (.A1(_02492_),
    .A2(_02493_),
    .B1(_02491_),
    .X(_02494_));
 sky130_fd_sc_hd__xor2_1 _08162_ (.A(_02485_),
    .B(_02486_),
    .X(_02495_));
 sky130_fd_sc_hd__a21o_1 _08163_ (.A1(_02494_),
    .A2(_02495_),
    .B1(_02488_),
    .X(_02496_));
 sky130_fd_sc_hd__xor2_1 _08164_ (.A(_02482_),
    .B(_02483_),
    .X(_02497_));
 sky130_fd_sc_hd__a21o_1 _08165_ (.A1(_02496_),
    .A2(_02497_),
    .B1(_02484_),
    .X(_02499_));
 sky130_fd_sc_hd__xor2_1 _08166_ (.A(_02479_),
    .B(_02480_),
    .X(_02500_));
 sky130_fd_sc_hd__a21o_1 _08167_ (.A1(_02499_),
    .A2(_02500_),
    .B1(_02481_),
    .X(_02501_));
 sky130_fd_sc_hd__xor2_1 _08168_ (.A(_02475_),
    .B(_02477_),
    .X(_02502_));
 sky130_fd_sc_hd__a21o_1 _08169_ (.A1(_02501_),
    .A2(_02502_),
    .B1(_02478_),
    .X(_02503_));
 sky130_fd_sc_hd__xor2_1 _08170_ (.A(_02472_),
    .B(_02473_),
    .X(_02504_));
 sky130_fd_sc_hd__a21o_1 _08171_ (.A1(_02503_),
    .A2(_02504_),
    .B1(_02474_),
    .X(_02505_));
 sky130_fd_sc_hd__xor2_1 _08172_ (.A(_02469_),
    .B(_02470_),
    .X(_02506_));
 sky130_fd_sc_hd__a21o_1 _08173_ (.A1(_02505_),
    .A2(_02506_),
    .B1(_02471_),
    .X(_02507_));
 sky130_fd_sc_hd__xor2_1 _08174_ (.A(_02466_),
    .B(_02467_),
    .X(_02508_));
 sky130_fd_sc_hd__a21o_1 _08175_ (.A1(_02507_),
    .A2(_02508_),
    .B1(_02468_),
    .X(_02510_));
 sky130_fd_sc_hd__xor2_1 _08176_ (.A(_02462_),
    .B(_02463_),
    .X(_02511_));
 sky130_fd_sc_hd__a21o_1 _08177_ (.A1(_02510_),
    .A2(_02511_),
    .B1(_02464_),
    .X(_02512_));
 sky130_fd_sc_hd__xor2_1 _08178_ (.A(_02459_),
    .B(_02460_),
    .X(_02513_));
 sky130_fd_sc_hd__a21o_1 _08179_ (.A1(_02512_),
    .A2(_02513_),
    .B1(_02461_),
    .X(_02514_));
 sky130_fd_sc_hd__xor2_1 _08180_ (.A(_02456_),
    .B(_02457_),
    .X(_02515_));
 sky130_fd_sc_hd__a21o_1 _08181_ (.A1(_02514_),
    .A2(_02515_),
    .B1(_02458_),
    .X(_02516_));
 sky130_fd_sc_hd__xor2_1 _08182_ (.A(_02452_),
    .B(_02453_),
    .X(_02517_));
 sky130_fd_sc_hd__a21o_1 _08183_ (.A1(_02516_),
    .A2(_02517_),
    .B1(_02455_),
    .X(_02518_));
 sky130_fd_sc_hd__xor2_1 _08184_ (.A(_02449_),
    .B(_02450_),
    .X(_02519_));
 sky130_fd_sc_hd__a21o_1 _08185_ (.A1(_02518_),
    .A2(_02519_),
    .B1(_02451_),
    .X(_02521_));
 sky130_fd_sc_hd__xor2_1 _08186_ (.A(_02446_),
    .B(_02447_),
    .X(_02522_));
 sky130_fd_sc_hd__a21o_1 _08187_ (.A1(_02521_),
    .A2(_02522_),
    .B1(_02448_),
    .X(_02523_));
 sky130_fd_sc_hd__xor2_1 _08188_ (.A(_02442_),
    .B(_02444_),
    .X(_02524_));
 sky130_fd_sc_hd__a21o_1 _08189_ (.A1(_02523_),
    .A2(_02524_),
    .B1(_02445_),
    .X(_02525_));
 sky130_fd_sc_hd__xor2_1 _08190_ (.A(_02439_),
    .B(_02440_),
    .X(_02526_));
 sky130_fd_sc_hd__a21oi_1 _08191_ (.A1(_02525_),
    .A2(_02526_),
    .B1(_02441_),
    .Y(_02527_));
 sky130_fd_sc_hd__nand2_1 _08192_ (.A(net41),
    .B(net25),
    .Y(_02528_));
 sky130_fd_sc_hd__and3_1 _08193_ (.A(_02340_),
    .B(_02430_),
    .C(_02528_),
    .X(_02529_));
 sky130_fd_sc_hd__and3_1 _08194_ (.A(net41),
    .B(net25),
    .C(_02431_),
    .X(_02530_));
 sky130_fd_sc_hd__nor2_1 _08195_ (.A(_02529_),
    .B(_02530_),
    .Y(_02532_));
 sky130_fd_sc_hd__a311o_1 _08196_ (.A1(net41),
    .A2(net24),
    .A3(_02435_),
    .B1(_02438_),
    .C1(_02532_),
    .X(_02533_));
 sky130_fd_sc_hd__nand2_1 _08197_ (.A(net42),
    .B(net24),
    .Y(_02534_));
 sky130_fd_sc_hd__xor2_1 _08198_ (.A(_02533_),
    .B(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__xnor2_1 _08199_ (.A(_02527_),
    .B(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__nand2_1 _08200_ (.A(net43),
    .B(net22),
    .Y(_02537_));
 sky130_fd_sc_hd__nor2_1 _08201_ (.A(_02536_),
    .B(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__xnor2_1 _08202_ (.A(_02525_),
    .B(_02526_),
    .Y(_02539_));
 sky130_fd_sc_hd__nand2_1 _08203_ (.A(net43),
    .B(net21),
    .Y(_02540_));
 sky130_fd_sc_hd__nor2_1 _08204_ (.A(_02539_),
    .B(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__xnor2_1 _08205_ (.A(_02523_),
    .B(_02524_),
    .Y(_02543_));
 sky130_fd_sc_hd__nand2_1 _08206_ (.A(net43),
    .B(net20),
    .Y(_02544_));
 sky130_fd_sc_hd__nor2_1 _08207_ (.A(_02543_),
    .B(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__xnor2_1 _08208_ (.A(_02521_),
    .B(_02522_),
    .Y(_02546_));
 sky130_fd_sc_hd__nand2_1 _08209_ (.A(net43),
    .B(net19),
    .Y(_02547_));
 sky130_fd_sc_hd__nor2_1 _08210_ (.A(_02546_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__xnor2_1 _08211_ (.A(_02518_),
    .B(_02519_),
    .Y(_02549_));
 sky130_fd_sc_hd__nand2_1 _08212_ (.A(net43),
    .B(net18),
    .Y(_02550_));
 sky130_fd_sc_hd__nor2_1 _08213_ (.A(_02549_),
    .B(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__xnor2_1 _08214_ (.A(_02516_),
    .B(_02517_),
    .Y(_02552_));
 sky130_fd_sc_hd__nand2_1 _08215_ (.A(net43),
    .B(net17),
    .Y(_02554_));
 sky130_fd_sc_hd__nor2_1 _08216_ (.A(_02552_),
    .B(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__xnor2_1 _08217_ (.A(_02514_),
    .B(_02515_),
    .Y(_02556_));
 sky130_fd_sc_hd__nand2_1 _08218_ (.A(net43),
    .B(net16),
    .Y(_02557_));
 sky130_fd_sc_hd__nor2_1 _08219_ (.A(_02556_),
    .B(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__xnor2_1 _08220_ (.A(_02512_),
    .B(_02513_),
    .Y(_02559_));
 sky130_fd_sc_hd__nand2_1 _08221_ (.A(net43),
    .B(net15),
    .Y(_02560_));
 sky130_fd_sc_hd__nor2_1 _08222_ (.A(_02559_),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__xnor2_1 _08223_ (.A(_02510_),
    .B(_02511_),
    .Y(_02562_));
 sky130_fd_sc_hd__nand2_1 _08224_ (.A(net43),
    .B(net14),
    .Y(_02563_));
 sky130_fd_sc_hd__nor2_1 _08225_ (.A(_02562_),
    .B(_02563_),
    .Y(_02565_));
 sky130_fd_sc_hd__xnor2_1 _08226_ (.A(_02507_),
    .B(_02508_),
    .Y(_02566_));
 sky130_fd_sc_hd__nand2_1 _08227_ (.A(net43),
    .B(net13),
    .Y(_02567_));
 sky130_fd_sc_hd__nor2_1 _08228_ (.A(_02566_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__xnor2_1 _08229_ (.A(_02505_),
    .B(_02506_),
    .Y(_02569_));
 sky130_fd_sc_hd__nand2_1 _08230_ (.A(net11),
    .B(net43),
    .Y(_02570_));
 sky130_fd_sc_hd__nor2_1 _08231_ (.A(_02569_),
    .B(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__xnor2_1 _08232_ (.A(_02503_),
    .B(_02504_),
    .Y(_02572_));
 sky130_fd_sc_hd__nand2_1 _08233_ (.A(net10),
    .B(net43),
    .Y(_02573_));
 sky130_fd_sc_hd__nor2_1 _08234_ (.A(_02572_),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__xnor2_1 _08235_ (.A(_02501_),
    .B(_02502_),
    .Y(_02576_));
 sky130_fd_sc_hd__nand2_1 _08236_ (.A(net9),
    .B(net43),
    .Y(_02577_));
 sky130_fd_sc_hd__nor2_1 _08237_ (.A(_02576_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__xnor2_1 _08238_ (.A(_02499_),
    .B(_02500_),
    .Y(_02579_));
 sky130_fd_sc_hd__nand2_1 _08239_ (.A(net8),
    .B(net43),
    .Y(_02580_));
 sky130_fd_sc_hd__nor2_1 _08240_ (.A(_02579_),
    .B(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__xnor2_1 _08241_ (.A(_02496_),
    .B(_02497_),
    .Y(_02582_));
 sky130_fd_sc_hd__nand2_1 _08242_ (.A(net7),
    .B(net43),
    .Y(_02583_));
 sky130_fd_sc_hd__nor2_1 _08243_ (.A(_02582_),
    .B(_02583_),
    .Y(_02584_));
 sky130_fd_sc_hd__xnor2_1 _08244_ (.A(_02494_),
    .B(_02495_),
    .Y(_02585_));
 sky130_fd_sc_hd__nand2_1 _08245_ (.A(net6),
    .B(net43),
    .Y(_02587_));
 sky130_fd_sc_hd__nor2_1 _08246_ (.A(_02585_),
    .B(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__xnor2_1 _08247_ (.A(_02492_),
    .B(_02493_),
    .Y(_02589_));
 sky130_fd_sc_hd__nand2_1 _08248_ (.A(net5),
    .B(net43),
    .Y(_02590_));
 sky130_fd_sc_hd__nor2_1 _08249_ (.A(_02589_),
    .B(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__a21o_1 _08250_ (.A1(_01492_),
    .A2(_01595_),
    .B1(_01594_),
    .X(_02592_));
 sky130_fd_sc_hd__xor2_1 _08251_ (.A(_02589_),
    .B(_02590_),
    .X(_02593_));
 sky130_fd_sc_hd__a21o_1 _08252_ (.A1(_02592_),
    .A2(_02593_),
    .B1(_02591_),
    .X(_02594_));
 sky130_fd_sc_hd__xor2_1 _08253_ (.A(_02585_),
    .B(_02587_),
    .X(_02595_));
 sky130_fd_sc_hd__a21o_1 _08254_ (.A1(_02594_),
    .A2(_02595_),
    .B1(_02588_),
    .X(_02596_));
 sky130_fd_sc_hd__xor2_1 _08255_ (.A(_02582_),
    .B(_02583_),
    .X(_02598_));
 sky130_fd_sc_hd__a21o_1 _08256_ (.A1(_02596_),
    .A2(_02598_),
    .B1(_02584_),
    .X(_02599_));
 sky130_fd_sc_hd__xor2_1 _08257_ (.A(_02579_),
    .B(_02580_),
    .X(_02600_));
 sky130_fd_sc_hd__a21o_1 _08258_ (.A1(_02599_),
    .A2(_02600_),
    .B1(_02581_),
    .X(_02601_));
 sky130_fd_sc_hd__xor2_1 _08259_ (.A(_02576_),
    .B(_02577_),
    .X(_02602_));
 sky130_fd_sc_hd__a21o_1 _08260_ (.A1(_02601_),
    .A2(_02602_),
    .B1(_02578_),
    .X(_02603_));
 sky130_fd_sc_hd__xor2_1 _08261_ (.A(_02572_),
    .B(_02573_),
    .X(_02604_));
 sky130_fd_sc_hd__a21o_1 _08262_ (.A1(_02603_),
    .A2(_02604_),
    .B1(_02574_),
    .X(_02605_));
 sky130_fd_sc_hd__xor2_1 _08263_ (.A(_02569_),
    .B(_02570_),
    .X(_02606_));
 sky130_fd_sc_hd__a21o_1 _08264_ (.A1(_02605_),
    .A2(_02606_),
    .B1(_02571_),
    .X(_02607_));
 sky130_fd_sc_hd__xor2_1 _08265_ (.A(_02566_),
    .B(_02567_),
    .X(_02609_));
 sky130_fd_sc_hd__a21o_1 _08266_ (.A1(_02607_),
    .A2(_02609_),
    .B1(_02568_),
    .X(_02610_));
 sky130_fd_sc_hd__xor2_1 _08267_ (.A(_02562_),
    .B(_02563_),
    .X(_02611_));
 sky130_fd_sc_hd__a21o_1 _08268_ (.A1(_02610_),
    .A2(_02611_),
    .B1(_02565_),
    .X(_02612_));
 sky130_fd_sc_hd__xor2_1 _08269_ (.A(_02559_),
    .B(_02560_),
    .X(_02613_));
 sky130_fd_sc_hd__a21o_1 _08270_ (.A1(_02612_),
    .A2(_02613_),
    .B1(_02561_),
    .X(_02614_));
 sky130_fd_sc_hd__xor2_1 _08271_ (.A(_02556_),
    .B(_02557_),
    .X(_02615_));
 sky130_fd_sc_hd__a21o_1 _08272_ (.A1(_02614_),
    .A2(_02615_),
    .B1(_02558_),
    .X(_02616_));
 sky130_fd_sc_hd__xor2_1 _08273_ (.A(_02552_),
    .B(_02554_),
    .X(_02617_));
 sky130_fd_sc_hd__a21o_1 _08274_ (.A1(_02616_),
    .A2(_02617_),
    .B1(_02555_),
    .X(_02618_));
 sky130_fd_sc_hd__xor2_1 _08275_ (.A(_02549_),
    .B(_02550_),
    .X(_02620_));
 sky130_fd_sc_hd__a21o_1 _08276_ (.A1(_02618_),
    .A2(_02620_),
    .B1(_02551_),
    .X(_02621_));
 sky130_fd_sc_hd__xor2_1 _08277_ (.A(_02546_),
    .B(_02547_),
    .X(_02622_));
 sky130_fd_sc_hd__a21o_1 _08278_ (.A1(_02621_),
    .A2(_02622_),
    .B1(_02548_),
    .X(_02623_));
 sky130_fd_sc_hd__xor2_1 _08279_ (.A(_02543_),
    .B(_02544_),
    .X(_02624_));
 sky130_fd_sc_hd__a21o_1 _08280_ (.A1(_02623_),
    .A2(_02624_),
    .B1(_02545_),
    .X(_02625_));
 sky130_fd_sc_hd__xor2_1 _08281_ (.A(_02539_),
    .B(_02540_),
    .X(_02626_));
 sky130_fd_sc_hd__a21o_1 _08282_ (.A1(_02625_),
    .A2(_02626_),
    .B1(_02541_),
    .X(_02627_));
 sky130_fd_sc_hd__xor2_1 _08283_ (.A(_02536_),
    .B(_02537_),
    .X(_02628_));
 sky130_fd_sc_hd__a21oi_1 _08284_ (.A1(_02627_),
    .A2(_02628_),
    .B1(_02538_),
    .Y(_02629_));
 sky130_fd_sc_hd__nand2_2 _08285_ (.A(net42),
    .B(net25),
    .Y(_02631_));
 sky130_fd_sc_hd__and2_1 _08286_ (.A(_02529_),
    .B(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__nor2_1 _08287_ (.A(_02529_),
    .B(_02631_),
    .Y(_02633_));
 sky130_fd_sc_hd__o22ai_1 _08288_ (.A1(_02527_),
    .A2(_02535_),
    .B1(_02632_),
    .B2(_02633_),
    .Y(_02634_));
 sky130_fd_sc_hd__a31o_1 _08289_ (.A1(net42),
    .A2(net24),
    .A3(_02533_),
    .B1(_02634_),
    .X(_02635_));
 sky130_fd_sc_hd__nand2_1 _08290_ (.A(net43),
    .B(net24),
    .Y(_02636_));
 sky130_fd_sc_hd__xor2_1 _08291_ (.A(_02635_),
    .B(_02636_),
    .X(_02637_));
 sky130_fd_sc_hd__nor2_1 _08292_ (.A(_02629_),
    .B(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__xnor2_1 _08293_ (.A(_02629_),
    .B(_02637_),
    .Y(_02639_));
 sky130_fd_sc_hd__nand2_1 _08294_ (.A(net45),
    .B(net22),
    .Y(_02640_));
 sky130_fd_sc_hd__nor2_1 _08295_ (.A(_02639_),
    .B(_02640_),
    .Y(_02642_));
 sky130_fd_sc_hd__xnor2_1 _08296_ (.A(_02627_),
    .B(_02628_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand2_1 _08297_ (.A(net45),
    .B(net21),
    .Y(_02644_));
 sky130_fd_sc_hd__nor2_1 _08298_ (.A(_02643_),
    .B(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__xnor2_1 _08299_ (.A(_02625_),
    .B(_02626_),
    .Y(_02646_));
 sky130_fd_sc_hd__nand2_1 _08300_ (.A(net45),
    .B(net20),
    .Y(_02647_));
 sky130_fd_sc_hd__nor2_1 _08301_ (.A(_02646_),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__xnor2_1 _08302_ (.A(_02623_),
    .B(_02624_),
    .Y(_02649_));
 sky130_fd_sc_hd__nand2_1 _08303_ (.A(net45),
    .B(net19),
    .Y(_02650_));
 sky130_fd_sc_hd__nor2_1 _08304_ (.A(_02649_),
    .B(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hd__xnor2_1 _08305_ (.A(_02621_),
    .B(_02622_),
    .Y(_02653_));
 sky130_fd_sc_hd__nand2_1 _08306_ (.A(net45),
    .B(net18),
    .Y(_02654_));
 sky130_fd_sc_hd__nor2_1 _08307_ (.A(_02653_),
    .B(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__xnor2_1 _08308_ (.A(_02618_),
    .B(_02620_),
    .Y(_02656_));
 sky130_fd_sc_hd__nand2_1 _08309_ (.A(net45),
    .B(net17),
    .Y(_02657_));
 sky130_fd_sc_hd__nor2_1 _08310_ (.A(_02656_),
    .B(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__xnor2_1 _08311_ (.A(_02616_),
    .B(_02617_),
    .Y(_02659_));
 sky130_fd_sc_hd__nand2_1 _08312_ (.A(net45),
    .B(net16),
    .Y(_02660_));
 sky130_fd_sc_hd__nor2_1 _08313_ (.A(_02659_),
    .B(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__xnor2_1 _08314_ (.A(_02614_),
    .B(_02615_),
    .Y(_02662_));
 sky130_fd_sc_hd__nand2_1 _08315_ (.A(net45),
    .B(net15),
    .Y(_02664_));
 sky130_fd_sc_hd__nor2_1 _08316_ (.A(_02662_),
    .B(_02664_),
    .Y(_02665_));
 sky130_fd_sc_hd__xnor2_1 _08317_ (.A(_02612_),
    .B(_02613_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand2_1 _08318_ (.A(net45),
    .B(net14),
    .Y(_02667_));
 sky130_fd_sc_hd__nor2_1 _08319_ (.A(_02666_),
    .B(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__xnor2_1 _08320_ (.A(_02610_),
    .B(_02611_),
    .Y(_02669_));
 sky130_fd_sc_hd__nand2_1 _08321_ (.A(net13),
    .B(net45),
    .Y(_02670_));
 sky130_fd_sc_hd__nor2_1 _08322_ (.A(_02669_),
    .B(_02670_),
    .Y(_02671_));
 sky130_fd_sc_hd__xnor2_1 _08323_ (.A(_02607_),
    .B(_02609_),
    .Y(_02672_));
 sky130_fd_sc_hd__nand2_1 _08324_ (.A(net11),
    .B(net45),
    .Y(_02673_));
 sky130_fd_sc_hd__nor2_1 _08325_ (.A(_02672_),
    .B(_02673_),
    .Y(_02675_));
 sky130_fd_sc_hd__xnor2_1 _08326_ (.A(_02605_),
    .B(_02606_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _08327_ (.A(net10),
    .B(net45),
    .Y(_02677_));
 sky130_fd_sc_hd__nor2_1 _08328_ (.A(_02676_),
    .B(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__xnor2_1 _08329_ (.A(_02603_),
    .B(_02604_),
    .Y(_02679_));
 sky130_fd_sc_hd__nand2_1 _08330_ (.A(net9),
    .B(net45),
    .Y(_02680_));
 sky130_fd_sc_hd__nor2_1 _08331_ (.A(_02679_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__xnor2_1 _08332_ (.A(_02601_),
    .B(_02602_),
    .Y(_02682_));
 sky130_fd_sc_hd__nand2_1 _08333_ (.A(net8),
    .B(net45),
    .Y(_02683_));
 sky130_fd_sc_hd__nor2_1 _08334_ (.A(_02682_),
    .B(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__xnor2_1 _08335_ (.A(_02599_),
    .B(_02600_),
    .Y(_02686_));
 sky130_fd_sc_hd__nand2_1 _08336_ (.A(net7),
    .B(net45),
    .Y(_02687_));
 sky130_fd_sc_hd__nor2_1 _08337_ (.A(_02686_),
    .B(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__xnor2_1 _08338_ (.A(_02596_),
    .B(_02598_),
    .Y(_02689_));
 sky130_fd_sc_hd__nand2_1 _08339_ (.A(net6),
    .B(net45),
    .Y(_02690_));
 sky130_fd_sc_hd__nor2_1 _08340_ (.A(_02689_),
    .B(_02690_),
    .Y(_02691_));
 sky130_fd_sc_hd__xnor2_1 _08341_ (.A(_02594_),
    .B(_02595_),
    .Y(_02692_));
 sky130_fd_sc_hd__nand2_1 _08342_ (.A(net5),
    .B(net45),
    .Y(_02693_));
 sky130_fd_sc_hd__nor2_1 _08343_ (.A(_02692_),
    .B(_02693_),
    .Y(_02694_));
 sky130_fd_sc_hd__xnor2_1 _08344_ (.A(_02592_),
    .B(_02593_),
    .Y(_02695_));
 sky130_fd_sc_hd__nand2_1 _08345_ (.A(net4),
    .B(net45),
    .Y(_02697_));
 sky130_fd_sc_hd__nor2_1 _08346_ (.A(_02695_),
    .B(_02697_),
    .Y(_02698_));
 sky130_fd_sc_hd__a21o_1 _08347_ (.A1(_01490_),
    .A2(_01599_),
    .B1(_01598_),
    .X(_02699_));
 sky130_fd_sc_hd__xor2_1 _08348_ (.A(_02695_),
    .B(_02697_),
    .X(_02700_));
 sky130_fd_sc_hd__a21o_1 _08349_ (.A1(_02699_),
    .A2(_02700_),
    .B1(_02698_),
    .X(_02701_));
 sky130_fd_sc_hd__xor2_1 _08350_ (.A(_02692_),
    .B(_02693_),
    .X(_02702_));
 sky130_fd_sc_hd__a21o_1 _08351_ (.A1(_02701_),
    .A2(_02702_),
    .B1(_02694_),
    .X(_02703_));
 sky130_fd_sc_hd__xor2_1 _08352_ (.A(_02689_),
    .B(_02690_),
    .X(_02704_));
 sky130_fd_sc_hd__a21o_1 _08353_ (.A1(_02703_),
    .A2(_02704_),
    .B1(_02691_),
    .X(_02705_));
 sky130_fd_sc_hd__xor2_1 _08354_ (.A(_02686_),
    .B(_02687_),
    .X(_02706_));
 sky130_fd_sc_hd__a21o_1 _08355_ (.A1(_02705_),
    .A2(_02706_),
    .B1(_02688_),
    .X(_02708_));
 sky130_fd_sc_hd__xor2_1 _08356_ (.A(_02682_),
    .B(_02683_),
    .X(_02709_));
 sky130_fd_sc_hd__a21o_1 _08357_ (.A1(_02708_),
    .A2(_02709_),
    .B1(_02684_),
    .X(_02710_));
 sky130_fd_sc_hd__xor2_1 _08358_ (.A(_02679_),
    .B(_02680_),
    .X(_02711_));
 sky130_fd_sc_hd__a21o_1 _08359_ (.A1(_02710_),
    .A2(_02711_),
    .B1(_02681_),
    .X(_02712_));
 sky130_fd_sc_hd__xor2_1 _08360_ (.A(_02676_),
    .B(_02677_),
    .X(_02713_));
 sky130_fd_sc_hd__a21o_1 _08361_ (.A1(_02712_),
    .A2(_02713_),
    .B1(_02678_),
    .X(_02714_));
 sky130_fd_sc_hd__xor2_1 _08362_ (.A(_02672_),
    .B(_02673_),
    .X(_02715_));
 sky130_fd_sc_hd__a21o_1 _08363_ (.A1(_02714_),
    .A2(_02715_),
    .B1(_02675_),
    .X(_02716_));
 sky130_fd_sc_hd__xor2_1 _08364_ (.A(_02669_),
    .B(_02670_),
    .X(_02717_));
 sky130_fd_sc_hd__a21o_1 _08365_ (.A1(_02716_),
    .A2(_02717_),
    .B1(_02671_),
    .X(_02719_));
 sky130_fd_sc_hd__xor2_1 _08366_ (.A(_02666_),
    .B(_02667_),
    .X(_02720_));
 sky130_fd_sc_hd__a21o_1 _08367_ (.A1(_02719_),
    .A2(_02720_),
    .B1(_02668_),
    .X(_02721_));
 sky130_fd_sc_hd__xor2_1 _08368_ (.A(_02662_),
    .B(_02664_),
    .X(_02722_));
 sky130_fd_sc_hd__a21o_1 _08369_ (.A1(_02721_),
    .A2(_02722_),
    .B1(_02665_),
    .X(_02723_));
 sky130_fd_sc_hd__xor2_1 _08370_ (.A(_02659_),
    .B(_02660_),
    .X(_02724_));
 sky130_fd_sc_hd__a21o_1 _08371_ (.A1(_02723_),
    .A2(_02724_),
    .B1(_02661_),
    .X(_02725_));
 sky130_fd_sc_hd__xor2_1 _08372_ (.A(_02656_),
    .B(_02657_),
    .X(_02726_));
 sky130_fd_sc_hd__a21o_1 _08373_ (.A1(_02725_),
    .A2(_02726_),
    .B1(_02658_),
    .X(_02727_));
 sky130_fd_sc_hd__xor2_1 _08374_ (.A(_02653_),
    .B(_02654_),
    .X(_02728_));
 sky130_fd_sc_hd__a21o_1 _08375_ (.A1(_02727_),
    .A2(_02728_),
    .B1(_02655_),
    .X(_02730_));
 sky130_fd_sc_hd__xor2_1 _08376_ (.A(_02649_),
    .B(_02650_),
    .X(_02731_));
 sky130_fd_sc_hd__a21o_1 _08377_ (.A1(_02730_),
    .A2(_02731_),
    .B1(_02651_),
    .X(_02732_));
 sky130_fd_sc_hd__xor2_1 _08378_ (.A(_02646_),
    .B(_02647_),
    .X(_02733_));
 sky130_fd_sc_hd__a21o_1 _08379_ (.A1(_02732_),
    .A2(_02733_),
    .B1(_02648_),
    .X(_02734_));
 sky130_fd_sc_hd__xor2_1 _08380_ (.A(_02643_),
    .B(_02644_),
    .X(_02735_));
 sky130_fd_sc_hd__a21o_1 _08381_ (.A1(_02734_),
    .A2(_02735_),
    .B1(_02645_),
    .X(_02736_));
 sky130_fd_sc_hd__xor2_1 _08382_ (.A(_02639_),
    .B(_02640_),
    .X(_02737_));
 sky130_fd_sc_hd__a21oi_1 _08383_ (.A1(_02736_),
    .A2(_02737_),
    .B1(_02642_),
    .Y(_02738_));
 sky130_fd_sc_hd__nand2_1 _08384_ (.A(net43),
    .B(net25),
    .Y(_02739_));
 sky130_fd_sc_hd__nand2_1 _08385_ (.A(_02632_),
    .B(_02739_),
    .Y(_02741_));
 sky130_fd_sc_hd__or2_1 _08386_ (.A(_02632_),
    .B(_02739_),
    .X(_02742_));
 sky130_fd_sc_hd__and2_1 _08387_ (.A(_02741_),
    .B(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__a311o_1 _08388_ (.A1(net43),
    .A2(net24),
    .A3(_02635_),
    .B1(_02638_),
    .C1(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__nand2_1 _08389_ (.A(net45),
    .B(net24),
    .Y(_02745_));
 sky130_fd_sc_hd__xor2_1 _08390_ (.A(_02744_),
    .B(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__xnor2_1 _08391_ (.A(_02738_),
    .B(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__nand2_1 _08392_ (.A(net46),
    .B(net22),
    .Y(_02748_));
 sky130_fd_sc_hd__nor2_1 _08393_ (.A(_02747_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__xnor2_1 _08394_ (.A(_02736_),
    .B(_02737_),
    .Y(_02750_));
 sky130_fd_sc_hd__nand2_1 _08395_ (.A(net46),
    .B(net21),
    .Y(_02752_));
 sky130_fd_sc_hd__nor2_1 _08396_ (.A(_02750_),
    .B(_02752_),
    .Y(_02753_));
 sky130_fd_sc_hd__xnor2_1 _08397_ (.A(_02734_),
    .B(_02735_),
    .Y(_02754_));
 sky130_fd_sc_hd__nand2_1 _08398_ (.A(net46),
    .B(net20),
    .Y(_02755_));
 sky130_fd_sc_hd__nor2_1 _08399_ (.A(_02754_),
    .B(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__xnor2_1 _08400_ (.A(_02732_),
    .B(_02733_),
    .Y(_02757_));
 sky130_fd_sc_hd__nand2_1 _08401_ (.A(net46),
    .B(net19),
    .Y(_02758_));
 sky130_fd_sc_hd__nor2_1 _08402_ (.A(_02757_),
    .B(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__xnor2_1 _08403_ (.A(_02730_),
    .B(_02731_),
    .Y(_02760_));
 sky130_fd_sc_hd__nand2_1 _08404_ (.A(net46),
    .B(net18),
    .Y(_02761_));
 sky130_fd_sc_hd__nor2_1 _08405_ (.A(_02760_),
    .B(_02761_),
    .Y(_02763_));
 sky130_fd_sc_hd__xnor2_1 _08406_ (.A(_02727_),
    .B(_02728_),
    .Y(_02764_));
 sky130_fd_sc_hd__nand2_1 _08407_ (.A(net46),
    .B(net17),
    .Y(_02765_));
 sky130_fd_sc_hd__nor2_1 _08408_ (.A(_02764_),
    .B(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__xnor2_1 _08409_ (.A(_02725_),
    .B(_02726_),
    .Y(_02767_));
 sky130_fd_sc_hd__nand2_1 _08410_ (.A(net46),
    .B(net16),
    .Y(_02768_));
 sky130_fd_sc_hd__nor2_1 _08411_ (.A(_02767_),
    .B(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__xnor2_1 _08412_ (.A(_02723_),
    .B(_02724_),
    .Y(_02770_));
 sky130_fd_sc_hd__nand2_1 _08413_ (.A(net46),
    .B(net15),
    .Y(_02771_));
 sky130_fd_sc_hd__nor2_1 _08414_ (.A(_02770_),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__xnor2_1 _08415_ (.A(_02721_),
    .B(_02722_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_1 _08416_ (.A(net14),
    .B(net46),
    .Y(_02775_));
 sky130_fd_sc_hd__nor2_1 _08417_ (.A(_02774_),
    .B(_02775_),
    .Y(_02776_));
 sky130_fd_sc_hd__xnor2_1 _08418_ (.A(_02719_),
    .B(_02720_),
    .Y(_02777_));
 sky130_fd_sc_hd__nand2_1 _08419_ (.A(net13),
    .B(net46),
    .Y(_02778_));
 sky130_fd_sc_hd__nor2_1 _08420_ (.A(_02777_),
    .B(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__xnor2_1 _08421_ (.A(_02716_),
    .B(_02717_),
    .Y(_02780_));
 sky130_fd_sc_hd__nand2_1 _08422_ (.A(net11),
    .B(net46),
    .Y(_02781_));
 sky130_fd_sc_hd__nor2_1 _08423_ (.A(_02780_),
    .B(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__xnor2_1 _08424_ (.A(_02714_),
    .B(_02715_),
    .Y(_02783_));
 sky130_fd_sc_hd__nand2_1 _08425_ (.A(net10),
    .B(net46),
    .Y(_02785_));
 sky130_fd_sc_hd__nor2_1 _08426_ (.A(_02783_),
    .B(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__xnor2_1 _08427_ (.A(_02712_),
    .B(_02713_),
    .Y(_02787_));
 sky130_fd_sc_hd__nand2_1 _08428_ (.A(net9),
    .B(net46),
    .Y(_02788_));
 sky130_fd_sc_hd__nor2_1 _08429_ (.A(_02787_),
    .B(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__xnor2_1 _08430_ (.A(_02710_),
    .B(_02711_),
    .Y(_02790_));
 sky130_fd_sc_hd__nand2_1 _08431_ (.A(net8),
    .B(net46),
    .Y(_02791_));
 sky130_fd_sc_hd__nor2_1 _08432_ (.A(_02790_),
    .B(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__xnor2_1 _08433_ (.A(_02708_),
    .B(_02709_),
    .Y(_02793_));
 sky130_fd_sc_hd__nand2_1 _08434_ (.A(net7),
    .B(net46),
    .Y(_02794_));
 sky130_fd_sc_hd__nor2_1 _08435_ (.A(_02793_),
    .B(_02794_),
    .Y(_02796_));
 sky130_fd_sc_hd__xnor2_1 _08436_ (.A(_02705_),
    .B(_02706_),
    .Y(_02797_));
 sky130_fd_sc_hd__nand2_1 _08437_ (.A(net6),
    .B(net46),
    .Y(_02798_));
 sky130_fd_sc_hd__nor2_1 _08438_ (.A(_02797_),
    .B(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__xnor2_1 _08439_ (.A(_02703_),
    .B(_02704_),
    .Y(_02800_));
 sky130_fd_sc_hd__nand2_1 _08440_ (.A(net5),
    .B(net46),
    .Y(_02801_));
 sky130_fd_sc_hd__nor2_1 _08441_ (.A(_02800_),
    .B(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__xnor2_1 _08442_ (.A(_02701_),
    .B(_02702_),
    .Y(_02803_));
 sky130_fd_sc_hd__nand2_1 _08443_ (.A(net4),
    .B(net46),
    .Y(_02804_));
 sky130_fd_sc_hd__nor2_1 _08444_ (.A(_02803_),
    .B(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__xnor2_1 _08445_ (.A(_02699_),
    .B(_02700_),
    .Y(_02807_));
 sky130_fd_sc_hd__nand2_1 _08446_ (.A(net3),
    .B(net46),
    .Y(_02808_));
 sky130_fd_sc_hd__nor2_1 _08447_ (.A(_02807_),
    .B(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__a21o_1 _08448_ (.A1(_01488_),
    .A2(_01602_),
    .B1(_01601_),
    .X(_02810_));
 sky130_fd_sc_hd__xor2_1 _08449_ (.A(_02807_),
    .B(_02808_),
    .X(_02811_));
 sky130_fd_sc_hd__a21o_1 _08450_ (.A1(_02810_),
    .A2(_02811_),
    .B1(_02809_),
    .X(_02812_));
 sky130_fd_sc_hd__xor2_1 _08451_ (.A(_02803_),
    .B(_02804_),
    .X(_02813_));
 sky130_fd_sc_hd__a21o_1 _08452_ (.A1(_02812_),
    .A2(_02813_),
    .B1(_02805_),
    .X(_02814_));
 sky130_fd_sc_hd__xor2_1 _08453_ (.A(_02800_),
    .B(_02801_),
    .X(_02815_));
 sky130_fd_sc_hd__a21o_1 _08454_ (.A1(_02814_),
    .A2(_02815_),
    .B1(_02802_),
    .X(_02816_));
 sky130_fd_sc_hd__xor2_1 _08455_ (.A(_02797_),
    .B(_02798_),
    .X(_02818_));
 sky130_fd_sc_hd__a21o_1 _08456_ (.A1(_02816_),
    .A2(_02818_),
    .B1(_02799_),
    .X(_02819_));
 sky130_fd_sc_hd__xor2_1 _08457_ (.A(_02793_),
    .B(_02794_),
    .X(_02820_));
 sky130_fd_sc_hd__a21o_1 _08458_ (.A1(_02819_),
    .A2(_02820_),
    .B1(_02796_),
    .X(_02821_));
 sky130_fd_sc_hd__xor2_1 _08459_ (.A(_02790_),
    .B(_02791_),
    .X(_02822_));
 sky130_fd_sc_hd__a21o_1 _08460_ (.A1(_02821_),
    .A2(_02822_),
    .B1(_02792_),
    .X(_02823_));
 sky130_fd_sc_hd__xor2_1 _08461_ (.A(_02787_),
    .B(_02788_),
    .X(_02824_));
 sky130_fd_sc_hd__a21o_1 _08462_ (.A1(_02823_),
    .A2(_02824_),
    .B1(_02789_),
    .X(_02825_));
 sky130_fd_sc_hd__xor2_1 _08463_ (.A(_02783_),
    .B(_02785_),
    .X(_02826_));
 sky130_fd_sc_hd__a21o_1 _08464_ (.A1(_02825_),
    .A2(_02826_),
    .B1(_02786_),
    .X(_02827_));
 sky130_fd_sc_hd__xor2_1 _08465_ (.A(_02780_),
    .B(_02781_),
    .X(_02829_));
 sky130_fd_sc_hd__a21o_1 _08466_ (.A1(_02827_),
    .A2(_02829_),
    .B1(_02782_),
    .X(_02830_));
 sky130_fd_sc_hd__xor2_1 _08467_ (.A(_02777_),
    .B(_02778_),
    .X(_02831_));
 sky130_fd_sc_hd__a21o_1 _08468_ (.A1(_02830_),
    .A2(_02831_),
    .B1(_02779_),
    .X(_02832_));
 sky130_fd_sc_hd__xor2_1 _08469_ (.A(_02774_),
    .B(_02775_),
    .X(_02833_));
 sky130_fd_sc_hd__a21o_1 _08470_ (.A1(_02832_),
    .A2(_02833_),
    .B1(_02776_),
    .X(_02834_));
 sky130_fd_sc_hd__xor2_1 _08471_ (.A(_02770_),
    .B(_02771_),
    .X(_02835_));
 sky130_fd_sc_hd__a21o_1 _08472_ (.A1(_02834_),
    .A2(_02835_),
    .B1(_02772_),
    .X(_02836_));
 sky130_fd_sc_hd__xor2_1 _08473_ (.A(_02767_),
    .B(_02768_),
    .X(_02837_));
 sky130_fd_sc_hd__a21o_1 _08474_ (.A1(_02836_),
    .A2(_02837_),
    .B1(_02769_),
    .X(_02838_));
 sky130_fd_sc_hd__xor2_1 _08475_ (.A(_02764_),
    .B(_02765_),
    .X(_02840_));
 sky130_fd_sc_hd__a21o_1 _08476_ (.A1(_02838_),
    .A2(_02840_),
    .B1(_02766_),
    .X(_02841_));
 sky130_fd_sc_hd__xor2_1 _08477_ (.A(_02760_),
    .B(_02761_),
    .X(_02842_));
 sky130_fd_sc_hd__a21o_1 _08478_ (.A1(_02841_),
    .A2(_02842_),
    .B1(_02763_),
    .X(_02843_));
 sky130_fd_sc_hd__xor2_1 _08479_ (.A(_02757_),
    .B(_02758_),
    .X(_02844_));
 sky130_fd_sc_hd__a21o_1 _08480_ (.A1(_02843_),
    .A2(_02844_),
    .B1(_02759_),
    .X(_02845_));
 sky130_fd_sc_hd__xor2_1 _08481_ (.A(_02754_),
    .B(_02755_),
    .X(_02846_));
 sky130_fd_sc_hd__a21o_1 _08482_ (.A1(_02845_),
    .A2(_02846_),
    .B1(_02756_),
    .X(_02847_));
 sky130_fd_sc_hd__xor2_1 _08483_ (.A(_02750_),
    .B(_02752_),
    .X(_02848_));
 sky130_fd_sc_hd__a21o_1 _08484_ (.A1(_02847_),
    .A2(_02848_),
    .B1(_02753_),
    .X(_02849_));
 sky130_fd_sc_hd__xor2_1 _08485_ (.A(_02747_),
    .B(_02748_),
    .X(_02851_));
 sky130_fd_sc_hd__a21oi_1 _08486_ (.A1(_02849_),
    .A2(_02851_),
    .B1(_02749_),
    .Y(_02852_));
 sky130_fd_sc_hd__nand2_1 _08487_ (.A(net45),
    .B(net25),
    .Y(_02853_));
 sky130_fd_sc_hd__nand2b_1 _08488_ (.A_N(_02741_),
    .B(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__a31o_1 _08489_ (.A1(_02529_),
    .A2(_02631_),
    .A3(_02739_),
    .B1(_02853_),
    .X(_02855_));
 sky130_fd_sc_hd__a2bb2o_1 _08490_ (.A1_N(_02738_),
    .A2_N(_02746_),
    .B1(_02854_),
    .B2(_02855_),
    .X(_02856_));
 sky130_fd_sc_hd__a31o_1 _08491_ (.A1(net45),
    .A2(net24),
    .A3(_02744_),
    .B1(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__nand2_1 _08492_ (.A(net46),
    .B(net24),
    .Y(_02858_));
 sky130_fd_sc_hd__and3_1 _08493_ (.A(net46),
    .B(net24),
    .C(_02857_),
    .X(_02859_));
 sky130_fd_sc_hd__xor2_1 _08494_ (.A(_02857_),
    .B(_02858_),
    .X(_02860_));
 sky130_fd_sc_hd__xnor2_1 _08495_ (.A(_02852_),
    .B(_02860_),
    .Y(_02862_));
 sky130_fd_sc_hd__nand2_1 _08496_ (.A(net47),
    .B(net22),
    .Y(_02863_));
 sky130_fd_sc_hd__nor2_1 _08497_ (.A(_02862_),
    .B(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__xnor2_1 _08498_ (.A(_02849_),
    .B(_02851_),
    .Y(_02865_));
 sky130_fd_sc_hd__nand2_1 _08499_ (.A(net47),
    .B(net21),
    .Y(_02866_));
 sky130_fd_sc_hd__nor2_1 _08500_ (.A(_02865_),
    .B(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__xnor2_1 _08501_ (.A(_02847_),
    .B(_02848_),
    .Y(_02868_));
 sky130_fd_sc_hd__nand2_1 _08502_ (.A(net47),
    .B(net20),
    .Y(_02869_));
 sky130_fd_sc_hd__nor2_1 _08503_ (.A(_02868_),
    .B(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__xnor2_1 _08504_ (.A(_02845_),
    .B(_02846_),
    .Y(_02871_));
 sky130_fd_sc_hd__nand2_1 _08505_ (.A(net47),
    .B(net19),
    .Y(_02873_));
 sky130_fd_sc_hd__nor2_1 _08506_ (.A(_02871_),
    .B(_02873_),
    .Y(_02874_));
 sky130_fd_sc_hd__xnor2_1 _08507_ (.A(_02843_),
    .B(_02844_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_1 _08508_ (.A(net47),
    .B(net18),
    .Y(_02876_));
 sky130_fd_sc_hd__nor2_1 _08509_ (.A(_02875_),
    .B(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__xnor2_1 _08510_ (.A(_02841_),
    .B(_02842_),
    .Y(_02878_));
 sky130_fd_sc_hd__nand2_1 _08511_ (.A(net47),
    .B(net17),
    .Y(_02879_));
 sky130_fd_sc_hd__nor2_1 _08512_ (.A(_02878_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__xnor2_1 _08513_ (.A(_02838_),
    .B(_02840_),
    .Y(_02881_));
 sky130_fd_sc_hd__nand2_1 _08514_ (.A(net47),
    .B(net16),
    .Y(_02882_));
 sky130_fd_sc_hd__nor2_1 _08515_ (.A(_02881_),
    .B(_02882_),
    .Y(_02884_));
 sky130_fd_sc_hd__xnor2_1 _08516_ (.A(_02836_),
    .B(_02837_),
    .Y(_02885_));
 sky130_fd_sc_hd__nand2_1 _08517_ (.A(net15),
    .B(net47),
    .Y(_02886_));
 sky130_fd_sc_hd__nor2_1 _08518_ (.A(_02885_),
    .B(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__xnor2_1 _08519_ (.A(_02834_),
    .B(_02835_),
    .Y(_02888_));
 sky130_fd_sc_hd__nand2_1 _08520_ (.A(net14),
    .B(net47),
    .Y(_02889_));
 sky130_fd_sc_hd__nor2_1 _08521_ (.A(_02888_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__xnor2_1 _08522_ (.A(_02832_),
    .B(_02833_),
    .Y(_02891_));
 sky130_fd_sc_hd__nand2_1 _08523_ (.A(net13),
    .B(net47),
    .Y(_02892_));
 sky130_fd_sc_hd__nor2_1 _08524_ (.A(_02891_),
    .B(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__xnor2_1 _08525_ (.A(_02830_),
    .B(_02831_),
    .Y(_02895_));
 sky130_fd_sc_hd__nand2_1 _08526_ (.A(net11),
    .B(net47),
    .Y(_02896_));
 sky130_fd_sc_hd__nor2_1 _08527_ (.A(_02895_),
    .B(_02896_),
    .Y(_02897_));
 sky130_fd_sc_hd__xnor2_1 _08528_ (.A(_02827_),
    .B(_02829_),
    .Y(_02898_));
 sky130_fd_sc_hd__nand2_1 _08529_ (.A(net10),
    .B(net47),
    .Y(_02899_));
 sky130_fd_sc_hd__nor2_1 _08530_ (.A(_02898_),
    .B(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__xnor2_1 _08531_ (.A(_02825_),
    .B(_02826_),
    .Y(_02901_));
 sky130_fd_sc_hd__nand2_1 _08532_ (.A(net9),
    .B(net47),
    .Y(_02902_));
 sky130_fd_sc_hd__nor2_1 _08533_ (.A(_02901_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__xnor2_1 _08534_ (.A(_02823_),
    .B(_02824_),
    .Y(_02904_));
 sky130_fd_sc_hd__nand2_1 _08535_ (.A(net8),
    .B(net47),
    .Y(_02906_));
 sky130_fd_sc_hd__nor2_1 _08536_ (.A(_02904_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__xnor2_1 _08537_ (.A(_02821_),
    .B(_02822_),
    .Y(_02908_));
 sky130_fd_sc_hd__nand2_1 _08538_ (.A(net7),
    .B(net47),
    .Y(_02909_));
 sky130_fd_sc_hd__nor2_1 _08539_ (.A(_02908_),
    .B(_02909_),
    .Y(_02910_));
 sky130_fd_sc_hd__xnor2_1 _08540_ (.A(_02819_),
    .B(_02820_),
    .Y(_02911_));
 sky130_fd_sc_hd__nand2_1 _08541_ (.A(net6),
    .B(net47),
    .Y(_02912_));
 sky130_fd_sc_hd__nor2_1 _08542_ (.A(_02911_),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__xnor2_1 _08543_ (.A(_02816_),
    .B(_02818_),
    .Y(_02914_));
 sky130_fd_sc_hd__nand2_1 _08544_ (.A(net5),
    .B(net47),
    .Y(_02915_));
 sky130_fd_sc_hd__nor2_1 _08545_ (.A(_02914_),
    .B(_02915_),
    .Y(_02917_));
 sky130_fd_sc_hd__xnor2_1 _08546_ (.A(_02814_),
    .B(_02815_),
    .Y(_02918_));
 sky130_fd_sc_hd__nand2_1 _08547_ (.A(net4),
    .B(net47),
    .Y(_02919_));
 sky130_fd_sc_hd__nor2_1 _08548_ (.A(_02918_),
    .B(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__xnor2_1 _08549_ (.A(_02812_),
    .B(_02813_),
    .Y(_02921_));
 sky130_fd_sc_hd__nand2_1 _08550_ (.A(net3),
    .B(net47),
    .Y(_02922_));
 sky130_fd_sc_hd__nor2_1 _08551_ (.A(_02921_),
    .B(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__xnor2_1 _08552_ (.A(_02810_),
    .B(_02811_),
    .Y(_02924_));
 sky130_fd_sc_hd__nand2_1 _08553_ (.A(net2),
    .B(net47),
    .Y(_02925_));
 sky130_fd_sc_hd__nor2_1 _08554_ (.A(_02924_),
    .B(_02925_),
    .Y(_02926_));
 sky130_fd_sc_hd__a21o_1 _08555_ (.A1(_01485_),
    .A2(_01605_),
    .B1(_01604_),
    .X(_02928_));
 sky130_fd_sc_hd__xor2_1 _08556_ (.A(_02924_),
    .B(_02925_),
    .X(_02929_));
 sky130_fd_sc_hd__a21o_1 _08557_ (.A1(_02928_),
    .A2(_02929_),
    .B1(_02926_),
    .X(_02930_));
 sky130_fd_sc_hd__xor2_1 _08558_ (.A(_02921_),
    .B(_02922_),
    .X(_02931_));
 sky130_fd_sc_hd__a21o_1 _08559_ (.A1(_02930_),
    .A2(_02931_),
    .B1(_02923_),
    .X(_02932_));
 sky130_fd_sc_hd__xor2_1 _08560_ (.A(_02918_),
    .B(_02919_),
    .X(_02933_));
 sky130_fd_sc_hd__a21o_1 _08561_ (.A1(_02932_),
    .A2(_02933_),
    .B1(_02920_),
    .X(_02934_));
 sky130_fd_sc_hd__xor2_1 _08562_ (.A(_02914_),
    .B(_02915_),
    .X(_02935_));
 sky130_fd_sc_hd__a21o_1 _08563_ (.A1(_02934_),
    .A2(_02935_),
    .B1(_02917_),
    .X(_02936_));
 sky130_fd_sc_hd__xor2_1 _08564_ (.A(_02911_),
    .B(_02912_),
    .X(_02937_));
 sky130_fd_sc_hd__a21o_1 _08565_ (.A1(_02936_),
    .A2(_02937_),
    .B1(_02913_),
    .X(_02939_));
 sky130_fd_sc_hd__xor2_1 _08566_ (.A(_02908_),
    .B(_02909_),
    .X(_02940_));
 sky130_fd_sc_hd__a21o_1 _08567_ (.A1(_02939_),
    .A2(_02940_),
    .B1(_02910_),
    .X(_02941_));
 sky130_fd_sc_hd__xor2_1 _08568_ (.A(_02904_),
    .B(_02906_),
    .X(_02942_));
 sky130_fd_sc_hd__a21o_1 _08569_ (.A1(_02941_),
    .A2(_02942_),
    .B1(_02907_),
    .X(_02943_));
 sky130_fd_sc_hd__xor2_1 _08570_ (.A(_02901_),
    .B(_02902_),
    .X(_02944_));
 sky130_fd_sc_hd__a21o_1 _08571_ (.A1(_02943_),
    .A2(_02944_),
    .B1(_02903_),
    .X(_02945_));
 sky130_fd_sc_hd__xor2_1 _08572_ (.A(_02898_),
    .B(_02899_),
    .X(_02946_));
 sky130_fd_sc_hd__a21o_1 _08573_ (.A1(_02945_),
    .A2(_02946_),
    .B1(_02900_),
    .X(_02947_));
 sky130_fd_sc_hd__xor2_1 _08574_ (.A(_02895_),
    .B(_02896_),
    .X(_02948_));
 sky130_fd_sc_hd__a21o_1 _08575_ (.A1(_02947_),
    .A2(_02948_),
    .B1(_02897_),
    .X(_02950_));
 sky130_fd_sc_hd__xor2_1 _08576_ (.A(_02891_),
    .B(_02892_),
    .X(_02951_));
 sky130_fd_sc_hd__a21o_1 _08577_ (.A1(_02950_),
    .A2(_02951_),
    .B1(_02893_),
    .X(_02952_));
 sky130_fd_sc_hd__xor2_1 _08578_ (.A(_02888_),
    .B(_02889_),
    .X(_02953_));
 sky130_fd_sc_hd__a21o_1 _08579_ (.A1(_02952_),
    .A2(_02953_),
    .B1(_02890_),
    .X(_02954_));
 sky130_fd_sc_hd__xor2_1 _08580_ (.A(_02885_),
    .B(_02886_),
    .X(_02955_));
 sky130_fd_sc_hd__a21o_1 _08581_ (.A1(_02954_),
    .A2(_02955_),
    .B1(_02887_),
    .X(_02956_));
 sky130_fd_sc_hd__xor2_1 _08582_ (.A(_02881_),
    .B(_02882_),
    .X(_02957_));
 sky130_fd_sc_hd__a21o_1 _08583_ (.A1(_02956_),
    .A2(_02957_),
    .B1(_02884_),
    .X(_02958_));
 sky130_fd_sc_hd__xor2_1 _08584_ (.A(_02878_),
    .B(_02879_),
    .X(_02959_));
 sky130_fd_sc_hd__a21o_1 _08585_ (.A1(_02958_),
    .A2(_02959_),
    .B1(_02880_),
    .X(_02961_));
 sky130_fd_sc_hd__xor2_1 _08586_ (.A(_02875_),
    .B(_02876_),
    .X(_02962_));
 sky130_fd_sc_hd__a21o_1 _08587_ (.A1(_02961_),
    .A2(_02962_),
    .B1(_02877_),
    .X(_02963_));
 sky130_fd_sc_hd__xor2_1 _08588_ (.A(_02871_),
    .B(_02873_),
    .X(_02964_));
 sky130_fd_sc_hd__a21o_1 _08589_ (.A1(_02963_),
    .A2(_02964_),
    .B1(_02874_),
    .X(_02965_));
 sky130_fd_sc_hd__xor2_1 _08590_ (.A(_02868_),
    .B(_02869_),
    .X(_02966_));
 sky130_fd_sc_hd__a21o_1 _08591_ (.A1(_02965_),
    .A2(_02966_),
    .B1(_02870_),
    .X(_02967_));
 sky130_fd_sc_hd__xor2_1 _08592_ (.A(_02865_),
    .B(_02866_),
    .X(_02968_));
 sky130_fd_sc_hd__a21o_1 _08593_ (.A1(_02967_),
    .A2(_02968_),
    .B1(_02867_),
    .X(_02969_));
 sky130_fd_sc_hd__xor2_1 _08594_ (.A(_02862_),
    .B(_02863_),
    .X(_02970_));
 sky130_fd_sc_hd__a21oi_1 _08595_ (.A1(_02969_),
    .A2(_02970_),
    .B1(_02864_),
    .Y(_02972_));
 sky130_fd_sc_hd__nand2_1 _08596_ (.A(net46),
    .B(net25),
    .Y(_02973_));
 sky130_fd_sc_hd__and2b_1 _08597_ (.A_N(_02854_),
    .B(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__and3_1 _08598_ (.A(net46),
    .B(net25),
    .C(_02854_),
    .X(_02975_));
 sky130_fd_sc_hd__o21ba_1 _08599_ (.A1(_02852_),
    .A2(_02860_),
    .B1_N(_02859_),
    .X(_02976_));
 sky130_fd_sc_hd__o21ai_1 _08600_ (.A1(_02974_),
    .A2(_02975_),
    .B1(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__nand2_1 _08601_ (.A(net47),
    .B(net24),
    .Y(_02978_));
 sky130_fd_sc_hd__xor2_1 _08602_ (.A(_02977_),
    .B(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__xnor2_1 _08603_ (.A(_02972_),
    .B(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__nand2_1 _08604_ (.A(net48),
    .B(net22),
    .Y(_02981_));
 sky130_fd_sc_hd__nor2_1 _08605_ (.A(_02980_),
    .B(_02981_),
    .Y(_02983_));
 sky130_fd_sc_hd__xnor2_1 _08606_ (.A(_02969_),
    .B(_02970_),
    .Y(_02984_));
 sky130_fd_sc_hd__nand2_1 _08607_ (.A(net48),
    .B(net21),
    .Y(_02985_));
 sky130_fd_sc_hd__nor2_1 _08608_ (.A(_02984_),
    .B(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hd__xnor2_1 _08609_ (.A(_02967_),
    .B(_02968_),
    .Y(_02987_));
 sky130_fd_sc_hd__nand2_1 _08610_ (.A(net48),
    .B(net20),
    .Y(_02988_));
 sky130_fd_sc_hd__nor2_1 _08611_ (.A(_02987_),
    .B(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__xnor2_1 _08612_ (.A(_02965_),
    .B(_02966_),
    .Y(_02990_));
 sky130_fd_sc_hd__nand2_1 _08613_ (.A(net48),
    .B(net19),
    .Y(_02991_));
 sky130_fd_sc_hd__nor2_1 _08614_ (.A(_02990_),
    .B(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__xnor2_1 _08615_ (.A(_02963_),
    .B(_02964_),
    .Y(_02994_));
 sky130_fd_sc_hd__nand2_1 _08616_ (.A(net48),
    .B(net18),
    .Y(_02995_));
 sky130_fd_sc_hd__nor2_1 _08617_ (.A(_02994_),
    .B(_02995_),
    .Y(_02996_));
 sky130_fd_sc_hd__xnor2_1 _08618_ (.A(_02961_),
    .B(_02962_),
    .Y(_02997_));
 sky130_fd_sc_hd__nand2_1 _08619_ (.A(net48),
    .B(net17),
    .Y(_02998_));
 sky130_fd_sc_hd__nor2_1 _08620_ (.A(_02997_),
    .B(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__xnor2_1 _08621_ (.A(_02958_),
    .B(_02959_),
    .Y(_03000_));
 sky130_fd_sc_hd__nand2_1 _08622_ (.A(net16),
    .B(net48),
    .Y(_03001_));
 sky130_fd_sc_hd__nor2_1 _08623_ (.A(_03000_),
    .B(_03001_),
    .Y(_03002_));
 sky130_fd_sc_hd__xnor2_1 _08624_ (.A(_02956_),
    .B(_02957_),
    .Y(_03003_));
 sky130_fd_sc_hd__nand2_1 _08625_ (.A(net15),
    .B(net48),
    .Y(_03005_));
 sky130_fd_sc_hd__nor2_1 _08626_ (.A(_03003_),
    .B(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__xnor2_1 _08627_ (.A(_02954_),
    .B(_02955_),
    .Y(_03007_));
 sky130_fd_sc_hd__nand2_1 _08628_ (.A(net14),
    .B(net48),
    .Y(_03008_));
 sky130_fd_sc_hd__nor2_1 _08629_ (.A(_03007_),
    .B(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__xnor2_1 _08630_ (.A(_02952_),
    .B(_02953_),
    .Y(_03010_));
 sky130_fd_sc_hd__nand2_1 _08631_ (.A(net13),
    .B(net48),
    .Y(_03011_));
 sky130_fd_sc_hd__nor2_1 _08632_ (.A(_03010_),
    .B(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__xnor2_1 _08633_ (.A(_02950_),
    .B(_02951_),
    .Y(_03013_));
 sky130_fd_sc_hd__nand2_1 _08634_ (.A(net11),
    .B(net48),
    .Y(_03014_));
 sky130_fd_sc_hd__nor2_1 _08635_ (.A(_03013_),
    .B(_03014_),
    .Y(_03016_));
 sky130_fd_sc_hd__xnor2_1 _08636_ (.A(_02947_),
    .B(_02948_),
    .Y(_03017_));
 sky130_fd_sc_hd__nand2_1 _08637_ (.A(net10),
    .B(net48),
    .Y(_03018_));
 sky130_fd_sc_hd__nor2_1 _08638_ (.A(_03017_),
    .B(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__xnor2_1 _08639_ (.A(_02945_),
    .B(_02946_),
    .Y(_03020_));
 sky130_fd_sc_hd__nand2_1 _08640_ (.A(net9),
    .B(net48),
    .Y(_03021_));
 sky130_fd_sc_hd__nor2_1 _08641_ (.A(_03020_),
    .B(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hd__xnor2_1 _08642_ (.A(_02943_),
    .B(_02944_),
    .Y(_03023_));
 sky130_fd_sc_hd__nand2_1 _08643_ (.A(net8),
    .B(net48),
    .Y(_03024_));
 sky130_fd_sc_hd__nor2_1 _08644_ (.A(_03023_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__xnor2_1 _08645_ (.A(_02941_),
    .B(_02942_),
    .Y(_03027_));
 sky130_fd_sc_hd__nand2_1 _08646_ (.A(net7),
    .B(net48),
    .Y(_03028_));
 sky130_fd_sc_hd__nor2_1 _08647_ (.A(_03027_),
    .B(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hd__xnor2_1 _08648_ (.A(_02939_),
    .B(_02940_),
    .Y(_03030_));
 sky130_fd_sc_hd__nand2_1 _08649_ (.A(net6),
    .B(net48),
    .Y(_03031_));
 sky130_fd_sc_hd__nor2_1 _08650_ (.A(_03030_),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__xnor2_1 _08651_ (.A(_02936_),
    .B(_02937_),
    .Y(_03033_));
 sky130_fd_sc_hd__nand2_1 _08652_ (.A(net5),
    .B(net48),
    .Y(_03034_));
 sky130_fd_sc_hd__nor2_1 _08653_ (.A(_03033_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__xnor2_1 _08654_ (.A(_02934_),
    .B(_02935_),
    .Y(_03036_));
 sky130_fd_sc_hd__nand2_1 _08655_ (.A(net4),
    .B(net48),
    .Y(_03038_));
 sky130_fd_sc_hd__nor2_1 _08656_ (.A(_03036_),
    .B(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__xnor2_1 _08657_ (.A(_02932_),
    .B(_02933_),
    .Y(_03040_));
 sky130_fd_sc_hd__nand2_1 _08658_ (.A(net3),
    .B(net48),
    .Y(_03041_));
 sky130_fd_sc_hd__nor2_1 _08659_ (.A(_03040_),
    .B(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__xnor2_1 _08660_ (.A(_02930_),
    .B(_02931_),
    .Y(_03043_));
 sky130_fd_sc_hd__nand2_1 _08661_ (.A(net2),
    .B(net48),
    .Y(_03044_));
 sky130_fd_sc_hd__nor2_1 _08662_ (.A(_03043_),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__xnor2_1 _08663_ (.A(_02928_),
    .B(_02929_),
    .Y(_03046_));
 sky130_fd_sc_hd__nand2_1 _08664_ (.A(net32),
    .B(net48),
    .Y(_03047_));
 sky130_fd_sc_hd__nor2_1 _08665_ (.A(_03046_),
    .B(_03047_),
    .Y(_03049_));
 sky130_fd_sc_hd__a21o_1 _08666_ (.A1(_01483_),
    .A2(_01609_),
    .B1(_01607_),
    .X(_03050_));
 sky130_fd_sc_hd__xor2_1 _08667_ (.A(_03046_),
    .B(_03047_),
    .X(_03051_));
 sky130_fd_sc_hd__a21o_1 _08668_ (.A1(_03050_),
    .A2(_03051_),
    .B1(_03049_),
    .X(_03052_));
 sky130_fd_sc_hd__xor2_1 _08669_ (.A(_03043_),
    .B(_03044_),
    .X(_03053_));
 sky130_fd_sc_hd__a21o_1 _08670_ (.A1(_03052_),
    .A2(_03053_),
    .B1(_03045_),
    .X(_03054_));
 sky130_fd_sc_hd__xor2_1 _08671_ (.A(_03040_),
    .B(_03041_),
    .X(_03055_));
 sky130_fd_sc_hd__a21o_1 _08672_ (.A1(_03054_),
    .A2(_03055_),
    .B1(_03042_),
    .X(_03056_));
 sky130_fd_sc_hd__xor2_1 _08673_ (.A(_03036_),
    .B(_03038_),
    .X(_03057_));
 sky130_fd_sc_hd__a21o_1 _08674_ (.A1(_03056_),
    .A2(_03057_),
    .B1(_03039_),
    .X(_03058_));
 sky130_fd_sc_hd__xor2_1 _08675_ (.A(_03033_),
    .B(_03034_),
    .X(_03060_));
 sky130_fd_sc_hd__a21o_1 _08676_ (.A1(_03058_),
    .A2(_03060_),
    .B1(_03035_),
    .X(_03061_));
 sky130_fd_sc_hd__xor2_1 _08677_ (.A(_03030_),
    .B(_03031_),
    .X(_03062_));
 sky130_fd_sc_hd__a21o_1 _08678_ (.A1(_03061_),
    .A2(_03062_),
    .B1(_03032_),
    .X(_03063_));
 sky130_fd_sc_hd__xor2_1 _08679_ (.A(_03027_),
    .B(_03028_),
    .X(_03064_));
 sky130_fd_sc_hd__a21o_1 _08680_ (.A1(_03063_),
    .A2(_03064_),
    .B1(_03029_),
    .X(_03065_));
 sky130_fd_sc_hd__xor2_1 _08681_ (.A(_03023_),
    .B(_03024_),
    .X(_03066_));
 sky130_fd_sc_hd__a21o_1 _08682_ (.A1(_03065_),
    .A2(_03066_),
    .B1(_03025_),
    .X(_03067_));
 sky130_fd_sc_hd__xor2_1 _08683_ (.A(_03020_),
    .B(_03021_),
    .X(_03068_));
 sky130_fd_sc_hd__a21o_1 _08684_ (.A1(_03067_),
    .A2(_03068_),
    .B1(_03022_),
    .X(_03069_));
 sky130_fd_sc_hd__xor2_1 _08685_ (.A(_03017_),
    .B(_03018_),
    .X(_03071_));
 sky130_fd_sc_hd__a21o_1 _08686_ (.A1(_03069_),
    .A2(_03071_),
    .B1(_03019_),
    .X(_03072_));
 sky130_fd_sc_hd__xor2_1 _08687_ (.A(_03013_),
    .B(_03014_),
    .X(_03073_));
 sky130_fd_sc_hd__a21o_1 _08688_ (.A1(_03072_),
    .A2(_03073_),
    .B1(_03016_),
    .X(_03074_));
 sky130_fd_sc_hd__xor2_1 _08689_ (.A(_03010_),
    .B(_03011_),
    .X(_03075_));
 sky130_fd_sc_hd__a21o_1 _08690_ (.A1(_03074_),
    .A2(_03075_),
    .B1(_03012_),
    .X(_03076_));
 sky130_fd_sc_hd__xor2_1 _08691_ (.A(_03007_),
    .B(_03008_),
    .X(_03077_));
 sky130_fd_sc_hd__a21o_1 _08692_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_03009_),
    .X(_03078_));
 sky130_fd_sc_hd__xor2_1 _08693_ (.A(_03003_),
    .B(_03005_),
    .X(_03079_));
 sky130_fd_sc_hd__a21o_1 _08694_ (.A1(_03078_),
    .A2(_03079_),
    .B1(_03006_),
    .X(_03080_));
 sky130_fd_sc_hd__xor2_1 _08695_ (.A(_03000_),
    .B(_03001_),
    .X(_03082_));
 sky130_fd_sc_hd__a21o_1 _08696_ (.A1(_03080_),
    .A2(_03082_),
    .B1(_03002_),
    .X(_03083_));
 sky130_fd_sc_hd__xor2_1 _08697_ (.A(_02997_),
    .B(_02998_),
    .X(_03084_));
 sky130_fd_sc_hd__a21o_1 _08698_ (.A1(_03083_),
    .A2(_03084_),
    .B1(_02999_),
    .X(_03085_));
 sky130_fd_sc_hd__xor2_1 _08699_ (.A(_02994_),
    .B(_02995_),
    .X(_03086_));
 sky130_fd_sc_hd__a21o_1 _08700_ (.A1(_03085_),
    .A2(_03086_),
    .B1(_02996_),
    .X(_03087_));
 sky130_fd_sc_hd__xor2_1 _08701_ (.A(_02990_),
    .B(_02991_),
    .X(_03088_));
 sky130_fd_sc_hd__a21o_1 _08702_ (.A1(_03087_),
    .A2(_03088_),
    .B1(_02992_),
    .X(_03089_));
 sky130_fd_sc_hd__xor2_1 _08703_ (.A(_02987_),
    .B(_02988_),
    .X(_03090_));
 sky130_fd_sc_hd__a21o_1 _08704_ (.A1(_03089_),
    .A2(_03090_),
    .B1(_02989_),
    .X(_03091_));
 sky130_fd_sc_hd__xor2_1 _08705_ (.A(_02984_),
    .B(_02985_),
    .X(_03093_));
 sky130_fd_sc_hd__a21o_1 _08706_ (.A1(_03091_),
    .A2(_03093_),
    .B1(_02986_),
    .X(_03094_));
 sky130_fd_sc_hd__xor2_1 _08707_ (.A(_02980_),
    .B(_02981_),
    .X(_03095_));
 sky130_fd_sc_hd__a21oi_1 _08708_ (.A1(_03094_),
    .A2(_03095_),
    .B1(_02983_),
    .Y(_03096_));
 sky130_fd_sc_hd__nand2_1 _08709_ (.A(net47),
    .B(net25),
    .Y(_03097_));
 sky130_fd_sc_hd__nand2_1 _08710_ (.A(_02974_),
    .B(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__or2_1 _08711_ (.A(_02974_),
    .B(_03097_),
    .X(_03099_));
 sky130_fd_sc_hd__a2bb2o_1 _08712_ (.A1_N(_02972_),
    .A2_N(_02979_),
    .B1(_03098_),
    .B2(_03099_),
    .X(_03100_));
 sky130_fd_sc_hd__a31o_1 _08713_ (.A1(net47),
    .A2(net24),
    .A3(_02977_),
    .B1(_03100_),
    .X(_03101_));
 sky130_fd_sc_hd__nand2_1 _08714_ (.A(net48),
    .B(net24),
    .Y(_03102_));
 sky130_fd_sc_hd__and3_1 _08715_ (.A(net48),
    .B(net24),
    .C(_03101_),
    .X(_03104_));
 sky130_fd_sc_hd__xor2_1 _08716_ (.A(_03101_),
    .B(_03102_),
    .X(_03105_));
 sky130_fd_sc_hd__xnor2_1 _08717_ (.A(_03096_),
    .B(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand2_1 _08718_ (.A(net49),
    .B(net22),
    .Y(_03107_));
 sky130_fd_sc_hd__nor2_1 _08719_ (.A(_03106_),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__xnor2_1 _08720_ (.A(_03094_),
    .B(_03095_),
    .Y(_03109_));
 sky130_fd_sc_hd__nand2_1 _08721_ (.A(net49),
    .B(net21),
    .Y(_03110_));
 sky130_fd_sc_hd__nor2_1 _08722_ (.A(_03109_),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__xnor2_1 _08723_ (.A(_03091_),
    .B(_03093_),
    .Y(_03112_));
 sky130_fd_sc_hd__nand2_1 _08724_ (.A(net49),
    .B(net20),
    .Y(_03113_));
 sky130_fd_sc_hd__nor2_1 _08725_ (.A(_03112_),
    .B(_03113_),
    .Y(_03115_));
 sky130_fd_sc_hd__xnor2_1 _08726_ (.A(_03089_),
    .B(_03090_),
    .Y(_03116_));
 sky130_fd_sc_hd__nand2_1 _08727_ (.A(net49),
    .B(net19),
    .Y(_03117_));
 sky130_fd_sc_hd__nor2_1 _08728_ (.A(_03116_),
    .B(_03117_),
    .Y(_03118_));
 sky130_fd_sc_hd__xnor2_1 _08729_ (.A(_03087_),
    .B(_03088_),
    .Y(_03119_));
 sky130_fd_sc_hd__nand2_1 _08730_ (.A(net49),
    .B(net18),
    .Y(_03120_));
 sky130_fd_sc_hd__nor2_1 _08731_ (.A(_03119_),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__xnor2_1 _08732_ (.A(_03085_),
    .B(_03086_),
    .Y(_03122_));
 sky130_fd_sc_hd__nand2_1 _08733_ (.A(net17),
    .B(net49),
    .Y(_03123_));
 sky130_fd_sc_hd__nor2_1 _08734_ (.A(_03122_),
    .B(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__xnor2_1 _08735_ (.A(_03083_),
    .B(_03084_),
    .Y(_03126_));
 sky130_fd_sc_hd__nand2_1 _08736_ (.A(net16),
    .B(net49),
    .Y(_03127_));
 sky130_fd_sc_hd__nor2_1 _08737_ (.A(_03126_),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__xnor2_1 _08738_ (.A(_03080_),
    .B(_03082_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand2_1 _08739_ (.A(net15),
    .B(net49),
    .Y(_03130_));
 sky130_fd_sc_hd__nor2_1 _08740_ (.A(_03129_),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__xnor2_1 _08741_ (.A(_03078_),
    .B(_03079_),
    .Y(_03132_));
 sky130_fd_sc_hd__nand2_1 _08742_ (.A(net14),
    .B(net49),
    .Y(_03133_));
 sky130_fd_sc_hd__nor2_1 _08743_ (.A(_03132_),
    .B(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__xnor2_1 _08744_ (.A(_03076_),
    .B(_03077_),
    .Y(_03135_));
 sky130_fd_sc_hd__nand2_1 _08745_ (.A(net13),
    .B(net49),
    .Y(_03137_));
 sky130_fd_sc_hd__nor2_1 _08746_ (.A(_03135_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__xnor2_1 _08747_ (.A(_03074_),
    .B(_03075_),
    .Y(_03139_));
 sky130_fd_sc_hd__nand2_1 _08748_ (.A(net11),
    .B(net49),
    .Y(_03140_));
 sky130_fd_sc_hd__nor2_1 _08749_ (.A(_03139_),
    .B(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__xnor2_1 _08750_ (.A(_03072_),
    .B(_03073_),
    .Y(_03142_));
 sky130_fd_sc_hd__nand2_1 _08751_ (.A(net10),
    .B(net49),
    .Y(_03143_));
 sky130_fd_sc_hd__nor2_1 _08752_ (.A(_03142_),
    .B(_03143_),
    .Y(_03144_));
 sky130_fd_sc_hd__xnor2_1 _08753_ (.A(_03069_),
    .B(_03071_),
    .Y(_03145_));
 sky130_fd_sc_hd__nand2_1 _08754_ (.A(net9),
    .B(net49),
    .Y(_03146_));
 sky130_fd_sc_hd__nor2_1 _08755_ (.A(_03145_),
    .B(_03146_),
    .Y(_03148_));
 sky130_fd_sc_hd__xnor2_1 _08756_ (.A(_03067_),
    .B(_03068_),
    .Y(_03149_));
 sky130_fd_sc_hd__nand2_1 _08757_ (.A(net8),
    .B(net49),
    .Y(_03150_));
 sky130_fd_sc_hd__nor2_1 _08758_ (.A(_03149_),
    .B(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__xnor2_1 _08759_ (.A(_03065_),
    .B(_03066_),
    .Y(_03152_));
 sky130_fd_sc_hd__nand2_1 _08760_ (.A(net7),
    .B(net49),
    .Y(_03153_));
 sky130_fd_sc_hd__nor2_1 _08761_ (.A(_03152_),
    .B(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__xnor2_1 _08762_ (.A(_03063_),
    .B(_03064_),
    .Y(_03155_));
 sky130_fd_sc_hd__nand2_1 _08763_ (.A(net6),
    .B(net49),
    .Y(_03156_));
 sky130_fd_sc_hd__nor2_1 _08764_ (.A(_03155_),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__xnor2_1 _08765_ (.A(_03061_),
    .B(_03062_),
    .Y(_03159_));
 sky130_fd_sc_hd__nand2_1 _08766_ (.A(net5),
    .B(net49),
    .Y(_03160_));
 sky130_fd_sc_hd__nor2_1 _08767_ (.A(_03159_),
    .B(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__xnor2_1 _08768_ (.A(_03058_),
    .B(_03060_),
    .Y(_03162_));
 sky130_fd_sc_hd__nand2_1 _08769_ (.A(net4),
    .B(net49),
    .Y(_03163_));
 sky130_fd_sc_hd__nor2_1 _08770_ (.A(_03162_),
    .B(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__xnor2_1 _08771_ (.A(_03056_),
    .B(_03057_),
    .Y(_03165_));
 sky130_fd_sc_hd__nand2_1 _08772_ (.A(net3),
    .B(net49),
    .Y(_03166_));
 sky130_fd_sc_hd__nor2_1 _08773_ (.A(_03165_),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__xnor2_1 _08774_ (.A(_03054_),
    .B(_03055_),
    .Y(_03168_));
 sky130_fd_sc_hd__nand2_1 _08775_ (.A(net2),
    .B(net49),
    .Y(_03170_));
 sky130_fd_sc_hd__nor2_1 _08776_ (.A(_03168_),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__xnor2_1 _08777_ (.A(_03052_),
    .B(_03053_),
    .Y(_03172_));
 sky130_fd_sc_hd__nand2_1 _08778_ (.A(net32),
    .B(net49),
    .Y(_03173_));
 sky130_fd_sc_hd__nor2_1 _08779_ (.A(_03172_),
    .B(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__xnor2_1 _08780_ (.A(_03050_),
    .B(_03051_),
    .Y(_03175_));
 sky130_fd_sc_hd__nand2_1 _08781_ (.A(net31),
    .B(net49),
    .Y(_03176_));
 sky130_fd_sc_hd__nor2_1 _08782_ (.A(_03175_),
    .B(_03176_),
    .Y(_03177_));
 sky130_fd_sc_hd__a21o_1 _08783_ (.A1(_01481_),
    .A2(_01612_),
    .B1(_01611_),
    .X(_03178_));
 sky130_fd_sc_hd__xor2_1 _08784_ (.A(_03175_),
    .B(_03176_),
    .X(_03179_));
 sky130_fd_sc_hd__a21o_1 _08785_ (.A1(_03178_),
    .A2(_03179_),
    .B1(_03177_),
    .X(_03181_));
 sky130_fd_sc_hd__xor2_1 _08786_ (.A(_03172_),
    .B(_03173_),
    .X(_03182_));
 sky130_fd_sc_hd__a21o_1 _08787_ (.A1(_03181_),
    .A2(_03182_),
    .B1(_03174_),
    .X(_03183_));
 sky130_fd_sc_hd__xor2_1 _08788_ (.A(_03168_),
    .B(_03170_),
    .X(_03184_));
 sky130_fd_sc_hd__a21o_1 _08789_ (.A1(_03183_),
    .A2(_03184_),
    .B1(_03171_),
    .X(_03185_));
 sky130_fd_sc_hd__xor2_1 _08790_ (.A(_03165_),
    .B(_03166_),
    .X(_03186_));
 sky130_fd_sc_hd__a21o_1 _08791_ (.A1(_03185_),
    .A2(_03186_),
    .B1(_03167_),
    .X(_03187_));
 sky130_fd_sc_hd__xor2_1 _08792_ (.A(_03162_),
    .B(_03163_),
    .X(_03188_));
 sky130_fd_sc_hd__a21o_1 _08793_ (.A1(_03187_),
    .A2(_03188_),
    .B1(_03164_),
    .X(_03189_));
 sky130_fd_sc_hd__xor2_1 _08794_ (.A(_03159_),
    .B(_03160_),
    .X(_03190_));
 sky130_fd_sc_hd__a21o_1 _08795_ (.A1(_03189_),
    .A2(_03190_),
    .B1(_03161_),
    .X(_03192_));
 sky130_fd_sc_hd__xor2_1 _08796_ (.A(_03155_),
    .B(_03156_),
    .X(_03193_));
 sky130_fd_sc_hd__a21o_1 _08797_ (.A1(_03192_),
    .A2(_03193_),
    .B1(_03157_),
    .X(_03194_));
 sky130_fd_sc_hd__xor2_1 _08798_ (.A(_03152_),
    .B(_03153_),
    .X(_03195_));
 sky130_fd_sc_hd__a21o_1 _08799_ (.A1(_03194_),
    .A2(_03195_),
    .B1(_03154_),
    .X(_03196_));
 sky130_fd_sc_hd__xor2_1 _08800_ (.A(_03149_),
    .B(_03150_),
    .X(_03197_));
 sky130_fd_sc_hd__a21o_1 _08801_ (.A1(_03196_),
    .A2(_03197_),
    .B1(_03151_),
    .X(_03198_));
 sky130_fd_sc_hd__xor2_1 _08802_ (.A(_03145_),
    .B(_03146_),
    .X(_03199_));
 sky130_fd_sc_hd__a21o_1 _08803_ (.A1(_03198_),
    .A2(_03199_),
    .B1(_03148_),
    .X(_03200_));
 sky130_fd_sc_hd__xor2_1 _08804_ (.A(_03142_),
    .B(_03143_),
    .X(_03201_));
 sky130_fd_sc_hd__a21o_1 _08805_ (.A1(_03200_),
    .A2(_03201_),
    .B1(_03144_),
    .X(_03203_));
 sky130_fd_sc_hd__xor2_1 _08806_ (.A(_03139_),
    .B(_03140_),
    .X(_03204_));
 sky130_fd_sc_hd__a21o_1 _08807_ (.A1(_03203_),
    .A2(_03204_),
    .B1(_03141_),
    .X(_03205_));
 sky130_fd_sc_hd__xor2_1 _08808_ (.A(_03135_),
    .B(_03137_),
    .X(_03206_));
 sky130_fd_sc_hd__a21o_1 _08809_ (.A1(_03205_),
    .A2(_03206_),
    .B1(_03138_),
    .X(_03207_));
 sky130_fd_sc_hd__xor2_1 _08810_ (.A(_03132_),
    .B(_03133_),
    .X(_03208_));
 sky130_fd_sc_hd__a21o_1 _08811_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03134_),
    .X(_03209_));
 sky130_fd_sc_hd__xor2_1 _08812_ (.A(_03129_),
    .B(_03130_),
    .X(_03210_));
 sky130_fd_sc_hd__a21o_1 _08813_ (.A1(_03209_),
    .A2(_03210_),
    .B1(_03131_),
    .X(_03211_));
 sky130_fd_sc_hd__xor2_1 _08814_ (.A(_03126_),
    .B(_03127_),
    .X(_03212_));
 sky130_fd_sc_hd__a21o_1 _08815_ (.A1(_03211_),
    .A2(_03212_),
    .B1(_03128_),
    .X(_03214_));
 sky130_fd_sc_hd__xor2_1 _08816_ (.A(_03122_),
    .B(_03123_),
    .X(_03215_));
 sky130_fd_sc_hd__a21o_1 _08817_ (.A1(_03214_),
    .A2(_03215_),
    .B1(_03124_),
    .X(_03216_));
 sky130_fd_sc_hd__xor2_1 _08818_ (.A(_03119_),
    .B(_03120_),
    .X(_03217_));
 sky130_fd_sc_hd__a21o_1 _08819_ (.A1(_03216_),
    .A2(_03217_),
    .B1(_03121_),
    .X(_03218_));
 sky130_fd_sc_hd__xor2_1 _08820_ (.A(_03116_),
    .B(_03117_),
    .X(_03219_));
 sky130_fd_sc_hd__a21o_1 _08821_ (.A1(_03218_),
    .A2(_03219_),
    .B1(_03118_),
    .X(_03220_));
 sky130_fd_sc_hd__xor2_1 _08822_ (.A(_03112_),
    .B(_03113_),
    .X(_03221_));
 sky130_fd_sc_hd__a21o_1 _08823_ (.A1(_03220_),
    .A2(_03221_),
    .B1(_03115_),
    .X(_03222_));
 sky130_fd_sc_hd__xor2_1 _08824_ (.A(_03109_),
    .B(_03110_),
    .X(_03223_));
 sky130_fd_sc_hd__a21o_1 _08825_ (.A1(_03222_),
    .A2(_03223_),
    .B1(_03111_),
    .X(_03225_));
 sky130_fd_sc_hd__xor2_1 _08826_ (.A(_03106_),
    .B(_03107_),
    .X(_03226_));
 sky130_fd_sc_hd__a21oi_1 _08827_ (.A1(_03225_),
    .A2(_03226_),
    .B1(_03108_),
    .Y(_03227_));
 sky130_fd_sc_hd__nand2_1 _08828_ (.A(net48),
    .B(net25),
    .Y(_03228_));
 sky130_fd_sc_hd__and3_1 _08829_ (.A(_02974_),
    .B(_03097_),
    .C(_03228_),
    .X(_03229_));
 sky130_fd_sc_hd__and3_1 _08830_ (.A(net48),
    .B(net25),
    .C(_03098_),
    .X(_03230_));
 sky130_fd_sc_hd__o21ba_1 _08831_ (.A1(_03096_),
    .A2(_03105_),
    .B1_N(_03104_),
    .X(_03231_));
 sky130_fd_sc_hd__o21ai_1 _08832_ (.A1(_03229_),
    .A2(_03230_),
    .B1(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__nand2_1 _08833_ (.A(net49),
    .B(net24),
    .Y(_03233_));
 sky130_fd_sc_hd__xor2_1 _08834_ (.A(_03232_),
    .B(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__xnor2_1 _08835_ (.A(_03227_),
    .B(_03234_),
    .Y(_03236_));
 sky130_fd_sc_hd__nand2_1 _08836_ (.A(net50),
    .B(net22),
    .Y(_03237_));
 sky130_fd_sc_hd__nor2_1 _08837_ (.A(_03236_),
    .B(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__xnor2_1 _08838_ (.A(_03225_),
    .B(_03226_),
    .Y(_03239_));
 sky130_fd_sc_hd__nand2_1 _08839_ (.A(net50),
    .B(net21),
    .Y(_03240_));
 sky130_fd_sc_hd__nor2_1 _08840_ (.A(_03239_),
    .B(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__xnor2_1 _08841_ (.A(_03222_),
    .B(_03223_),
    .Y(_03242_));
 sky130_fd_sc_hd__nand2_1 _08842_ (.A(net50),
    .B(net20),
    .Y(_03243_));
 sky130_fd_sc_hd__nor2_1 _08843_ (.A(_03242_),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__xnor2_1 _08844_ (.A(_03220_),
    .B(_03221_),
    .Y(_03245_));
 sky130_fd_sc_hd__nand2_1 _08845_ (.A(net50),
    .B(net19),
    .Y(_03247_));
 sky130_fd_sc_hd__nor2_1 _08846_ (.A(_03245_),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__xnor2_1 _08847_ (.A(_03218_),
    .B(_03219_),
    .Y(_03249_));
 sky130_fd_sc_hd__nand2_1 _08848_ (.A(net18),
    .B(net50),
    .Y(_03250_));
 sky130_fd_sc_hd__nor2_1 _08849_ (.A(_03249_),
    .B(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__xnor2_1 _08850_ (.A(_03216_),
    .B(_03217_),
    .Y(_03252_));
 sky130_fd_sc_hd__nand2_1 _08851_ (.A(net17),
    .B(net50),
    .Y(_03253_));
 sky130_fd_sc_hd__nor2_1 _08852_ (.A(_03252_),
    .B(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__xnor2_1 _08853_ (.A(_03214_),
    .B(_03215_),
    .Y(_03255_));
 sky130_fd_sc_hd__nand2_1 _08854_ (.A(net16),
    .B(net50),
    .Y(_03256_));
 sky130_fd_sc_hd__nor2_1 _08855_ (.A(_03255_),
    .B(_03256_),
    .Y(_03258_));
 sky130_fd_sc_hd__xnor2_1 _08856_ (.A(_03211_),
    .B(_03212_),
    .Y(_03259_));
 sky130_fd_sc_hd__nand2_1 _08857_ (.A(net15),
    .B(net50),
    .Y(_03260_));
 sky130_fd_sc_hd__nor2_1 _08858_ (.A(_03259_),
    .B(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__xnor2_1 _08859_ (.A(_03209_),
    .B(_03210_),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _08860_ (.A(net14),
    .B(net50),
    .Y(_03263_));
 sky130_fd_sc_hd__nor2_1 _08861_ (.A(_03262_),
    .B(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__xnor2_1 _08862_ (.A(_03207_),
    .B(_03208_),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2_1 _08863_ (.A(net13),
    .B(net50),
    .Y(_03266_));
 sky130_fd_sc_hd__nor2_1 _08864_ (.A(_03265_),
    .B(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__xnor2_1 _08865_ (.A(_03205_),
    .B(_03206_),
    .Y(_03269_));
 sky130_fd_sc_hd__nand2_1 _08866_ (.A(net11),
    .B(net50),
    .Y(_03270_));
 sky130_fd_sc_hd__nor2_1 _08867_ (.A(_03269_),
    .B(_03270_),
    .Y(_03271_));
 sky130_fd_sc_hd__xnor2_1 _08868_ (.A(_03203_),
    .B(_03204_),
    .Y(_03272_));
 sky130_fd_sc_hd__nand2_1 _08869_ (.A(net10),
    .B(net50),
    .Y(_03273_));
 sky130_fd_sc_hd__nor2_1 _08870_ (.A(_03272_),
    .B(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__xnor2_1 _08871_ (.A(_03200_),
    .B(_03201_),
    .Y(_03275_));
 sky130_fd_sc_hd__nand2_1 _08872_ (.A(net9),
    .B(net50),
    .Y(_03276_));
 sky130_fd_sc_hd__nor2_1 _08873_ (.A(_03275_),
    .B(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__xnor2_1 _08874_ (.A(_03198_),
    .B(_03199_),
    .Y(_03278_));
 sky130_fd_sc_hd__nand2_1 _08875_ (.A(net8),
    .B(net50),
    .Y(_03280_));
 sky130_fd_sc_hd__nor2_1 _08876_ (.A(_03278_),
    .B(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__xnor2_1 _08877_ (.A(_03196_),
    .B(_03197_),
    .Y(_03282_));
 sky130_fd_sc_hd__nand2_1 _08878_ (.A(net7),
    .B(net50),
    .Y(_03283_));
 sky130_fd_sc_hd__nor2_1 _08879_ (.A(_03282_),
    .B(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__xnor2_1 _08880_ (.A(_03194_),
    .B(_03195_),
    .Y(_03285_));
 sky130_fd_sc_hd__nand2_1 _08881_ (.A(net6),
    .B(net50),
    .Y(_03286_));
 sky130_fd_sc_hd__nor2_1 _08882_ (.A(_03285_),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__xnor2_1 _08883_ (.A(_03192_),
    .B(_03193_),
    .Y(_03288_));
 sky130_fd_sc_hd__nand2_1 _08884_ (.A(net5),
    .B(net50),
    .Y(_03289_));
 sky130_fd_sc_hd__nor2_1 _08885_ (.A(_03288_),
    .B(_03289_),
    .Y(_03291_));
 sky130_fd_sc_hd__xnor2_1 _08886_ (.A(_03189_),
    .B(_03190_),
    .Y(_03292_));
 sky130_fd_sc_hd__nand2_1 _08887_ (.A(net4),
    .B(net50),
    .Y(_03293_));
 sky130_fd_sc_hd__nor2_1 _08888_ (.A(_03292_),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__xnor2_1 _08889_ (.A(_03187_),
    .B(_03188_),
    .Y(_03295_));
 sky130_fd_sc_hd__nand2_1 _08890_ (.A(net3),
    .B(net50),
    .Y(_03296_));
 sky130_fd_sc_hd__nor2_1 _08891_ (.A(_03295_),
    .B(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__xnor2_1 _08892_ (.A(_03185_),
    .B(_03186_),
    .Y(_03298_));
 sky130_fd_sc_hd__nand2_1 _08893_ (.A(net2),
    .B(net50),
    .Y(_03299_));
 sky130_fd_sc_hd__nor2_1 _08894_ (.A(_03298_),
    .B(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__xnor2_1 _08895_ (.A(_03183_),
    .B(_03184_),
    .Y(_03302_));
 sky130_fd_sc_hd__nand2_1 _08896_ (.A(net32),
    .B(net50),
    .Y(_03303_));
 sky130_fd_sc_hd__nor2_1 _08897_ (.A(_03302_),
    .B(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__xnor2_1 _08898_ (.A(_03181_),
    .B(_03182_),
    .Y(_03305_));
 sky130_fd_sc_hd__nand2_1 _08899_ (.A(net31),
    .B(net50),
    .Y(_03306_));
 sky130_fd_sc_hd__nor2_1 _08900_ (.A(_03305_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__xnor2_1 _08901_ (.A(_03178_),
    .B(_03179_),
    .Y(_03308_));
 sky130_fd_sc_hd__nand2_1 _08902_ (.A(net30),
    .B(net50),
    .Y(_03309_));
 sky130_fd_sc_hd__nor2_1 _08903_ (.A(_03308_),
    .B(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__a21o_1 _08904_ (.A1(_01479_),
    .A2(_01615_),
    .B1(_01614_),
    .X(_03311_));
 sky130_fd_sc_hd__xor2_1 _08905_ (.A(_03308_),
    .B(_03309_),
    .X(_03313_));
 sky130_fd_sc_hd__a21o_1 _08906_ (.A1(_03311_),
    .A2(_03313_),
    .B1(_03310_),
    .X(_03314_));
 sky130_fd_sc_hd__xor2_1 _08907_ (.A(_03305_),
    .B(_03306_),
    .X(_03315_));
 sky130_fd_sc_hd__a21o_1 _08908_ (.A1(_03314_),
    .A2(_03315_),
    .B1(_03307_),
    .X(_03316_));
 sky130_fd_sc_hd__xor2_1 _08909_ (.A(_03302_),
    .B(_03303_),
    .X(_03317_));
 sky130_fd_sc_hd__a21o_1 _08910_ (.A1(_03316_),
    .A2(_03317_),
    .B1(_03304_),
    .X(_03318_));
 sky130_fd_sc_hd__xor2_1 _08911_ (.A(_03298_),
    .B(_03299_),
    .X(_03319_));
 sky130_fd_sc_hd__a21o_1 _08912_ (.A1(_03318_),
    .A2(_03319_),
    .B1(_03300_),
    .X(_03320_));
 sky130_fd_sc_hd__xor2_1 _08913_ (.A(_03295_),
    .B(_03296_),
    .X(_03321_));
 sky130_fd_sc_hd__a21o_1 _08914_ (.A1(_03320_),
    .A2(_03321_),
    .B1(_03297_),
    .X(_03322_));
 sky130_fd_sc_hd__xor2_1 _08915_ (.A(_03292_),
    .B(_03293_),
    .X(_03324_));
 sky130_fd_sc_hd__a21o_1 _08916_ (.A1(_03322_),
    .A2(_03324_),
    .B1(_03294_),
    .X(_03325_));
 sky130_fd_sc_hd__xor2_1 _08917_ (.A(_03288_),
    .B(_03289_),
    .X(_03326_));
 sky130_fd_sc_hd__a21o_1 _08918_ (.A1(_03325_),
    .A2(_03326_),
    .B1(_03291_),
    .X(_03327_));
 sky130_fd_sc_hd__xor2_1 _08919_ (.A(_03285_),
    .B(_03286_),
    .X(_03328_));
 sky130_fd_sc_hd__a21o_1 _08920_ (.A1(_03327_),
    .A2(_03328_),
    .B1(_03287_),
    .X(_03329_));
 sky130_fd_sc_hd__xor2_1 _08921_ (.A(_03282_),
    .B(_03283_),
    .X(_03330_));
 sky130_fd_sc_hd__a21o_1 _08922_ (.A1(_03329_),
    .A2(_03330_),
    .B1(_03284_),
    .X(_03331_));
 sky130_fd_sc_hd__xor2_1 _08923_ (.A(_03278_),
    .B(_03280_),
    .X(_03332_));
 sky130_fd_sc_hd__a21o_1 _08924_ (.A1(_03331_),
    .A2(_03332_),
    .B1(_03281_),
    .X(_03333_));
 sky130_fd_sc_hd__xor2_1 _08925_ (.A(_03275_),
    .B(_03276_),
    .X(_03335_));
 sky130_fd_sc_hd__a21o_1 _08926_ (.A1(_03333_),
    .A2(_03335_),
    .B1(_03277_),
    .X(_03336_));
 sky130_fd_sc_hd__xor2_1 _08927_ (.A(_03272_),
    .B(_03273_),
    .X(_03337_));
 sky130_fd_sc_hd__a21o_1 _08928_ (.A1(_03336_),
    .A2(_03337_),
    .B1(_03274_),
    .X(_03338_));
 sky130_fd_sc_hd__xor2_1 _08929_ (.A(_03269_),
    .B(_03270_),
    .X(_03339_));
 sky130_fd_sc_hd__a21o_1 _08930_ (.A1(_03338_),
    .A2(_03339_),
    .B1(_03271_),
    .X(_03340_));
 sky130_fd_sc_hd__xor2_1 _08931_ (.A(_03265_),
    .B(_03266_),
    .X(_03341_));
 sky130_fd_sc_hd__a21o_1 _08932_ (.A1(_03340_),
    .A2(_03341_),
    .B1(_03267_),
    .X(_03342_));
 sky130_fd_sc_hd__xor2_1 _08933_ (.A(_03262_),
    .B(_03263_),
    .X(_03343_));
 sky130_fd_sc_hd__a21o_1 _08934_ (.A1(_03342_),
    .A2(_03343_),
    .B1(_03264_),
    .X(_03344_));
 sky130_fd_sc_hd__xor2_1 _08935_ (.A(_03259_),
    .B(_03260_),
    .X(_03346_));
 sky130_fd_sc_hd__a21o_1 _08936_ (.A1(_03344_),
    .A2(_03346_),
    .B1(_03261_),
    .X(_03347_));
 sky130_fd_sc_hd__xor2_1 _08937_ (.A(_03255_),
    .B(_03256_),
    .X(_03348_));
 sky130_fd_sc_hd__a21o_1 _08938_ (.A1(_03347_),
    .A2(_03348_),
    .B1(_03258_),
    .X(_03349_));
 sky130_fd_sc_hd__xor2_1 _08939_ (.A(_03252_),
    .B(_03253_),
    .X(_03350_));
 sky130_fd_sc_hd__a21o_1 _08940_ (.A1(_03349_),
    .A2(_03350_),
    .B1(_03254_),
    .X(_03351_));
 sky130_fd_sc_hd__xor2_1 _08941_ (.A(_03249_),
    .B(_03250_),
    .X(_03352_));
 sky130_fd_sc_hd__a21o_1 _08942_ (.A1(_03351_),
    .A2(_03352_),
    .B1(_03251_),
    .X(_03353_));
 sky130_fd_sc_hd__xor2_1 _08943_ (.A(_03245_),
    .B(_03247_),
    .X(_03354_));
 sky130_fd_sc_hd__a21o_1 _08944_ (.A1(_03353_),
    .A2(_03354_),
    .B1(_03248_),
    .X(_03355_));
 sky130_fd_sc_hd__xor2_1 _08945_ (.A(_03242_),
    .B(_03243_),
    .X(_03357_));
 sky130_fd_sc_hd__a21o_1 _08946_ (.A1(_03355_),
    .A2(_03357_),
    .B1(_03244_),
    .X(_03358_));
 sky130_fd_sc_hd__xor2_1 _08947_ (.A(_03239_),
    .B(_03240_),
    .X(_03359_));
 sky130_fd_sc_hd__a21o_1 _08948_ (.A1(_03358_),
    .A2(_03359_),
    .B1(_03241_),
    .X(_03360_));
 sky130_fd_sc_hd__xor2_1 _08949_ (.A(_03236_),
    .B(_03237_),
    .X(_03361_));
 sky130_fd_sc_hd__a21oi_1 _08950_ (.A1(_03360_),
    .A2(_03361_),
    .B1(_03238_),
    .Y(_03362_));
 sky130_fd_sc_hd__nand2_1 _08951_ (.A(net49),
    .B(net25),
    .Y(_03363_));
 sky130_fd_sc_hd__and2_1 _08952_ (.A(_03229_),
    .B(_03363_),
    .X(_03364_));
 sky130_fd_sc_hd__nor2_1 _08953_ (.A(_03229_),
    .B(_03363_),
    .Y(_03365_));
 sky130_fd_sc_hd__o22ai_1 _08954_ (.A1(_03227_),
    .A2(_03234_),
    .B1(_03364_),
    .B2(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__a31o_1 _08955_ (.A1(net49),
    .A2(net24),
    .A3(_03232_),
    .B1(_03366_),
    .X(_03368_));
 sky130_fd_sc_hd__nand2_1 _08956_ (.A(net50),
    .B(net24),
    .Y(_03369_));
 sky130_fd_sc_hd__xor2_1 _08957_ (.A(_03368_),
    .B(_03369_),
    .X(_03370_));
 sky130_fd_sc_hd__xnor2_1 _08958_ (.A(_03362_),
    .B(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand2_1 _08959_ (.A(net51),
    .B(net22),
    .Y(_03372_));
 sky130_fd_sc_hd__nor2_1 _08960_ (.A(_03371_),
    .B(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__xnor2_1 _08961_ (.A(_03360_),
    .B(_03361_),
    .Y(_03374_));
 sky130_fd_sc_hd__nand2_1 _08962_ (.A(net51),
    .B(net21),
    .Y(_03375_));
 sky130_fd_sc_hd__nor2_1 _08963_ (.A(_03374_),
    .B(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__xnor2_1 _08964_ (.A(_03358_),
    .B(_03359_),
    .Y(_03377_));
 sky130_fd_sc_hd__nand2_1 _08965_ (.A(net51),
    .B(net20),
    .Y(_03379_));
 sky130_fd_sc_hd__nor2_1 _08966_ (.A(_03377_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__xnor2_1 _08967_ (.A(_03355_),
    .B(_03357_),
    .Y(_03381_));
 sky130_fd_sc_hd__nand2_1 _08968_ (.A(net19),
    .B(net51),
    .Y(_03382_));
 sky130_fd_sc_hd__nor2_1 _08969_ (.A(_03381_),
    .B(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__xnor2_1 _08970_ (.A(_03353_),
    .B(_03354_),
    .Y(_03384_));
 sky130_fd_sc_hd__nand2_1 _08971_ (.A(net18),
    .B(net51),
    .Y(_03385_));
 sky130_fd_sc_hd__nor2_1 _08972_ (.A(_03384_),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__xnor2_1 _08973_ (.A(_03351_),
    .B(_03352_),
    .Y(_03387_));
 sky130_fd_sc_hd__nand2_1 _08974_ (.A(net17),
    .B(net51),
    .Y(_03388_));
 sky130_fd_sc_hd__nor2_1 _08975_ (.A(_03387_),
    .B(_03388_),
    .Y(_03390_));
 sky130_fd_sc_hd__xnor2_1 _08976_ (.A(_03349_),
    .B(_03350_),
    .Y(_03391_));
 sky130_fd_sc_hd__nand2_1 _08977_ (.A(net16),
    .B(net51),
    .Y(_03392_));
 sky130_fd_sc_hd__nor2_1 _08978_ (.A(_03391_),
    .B(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__xnor2_1 _08979_ (.A(_03347_),
    .B(_03348_),
    .Y(_03394_));
 sky130_fd_sc_hd__nand2_1 _08980_ (.A(net15),
    .B(net51),
    .Y(_03395_));
 sky130_fd_sc_hd__nor2_1 _08981_ (.A(_03394_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__xnor2_1 _08982_ (.A(_03344_),
    .B(_03346_),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_1 _08983_ (.A(net14),
    .B(net51),
    .Y(_03398_));
 sky130_fd_sc_hd__nor2_1 _08984_ (.A(_03397_),
    .B(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__xnor2_1 _08985_ (.A(_03342_),
    .B(_03343_),
    .Y(_03401_));
 sky130_fd_sc_hd__nand2_1 _08986_ (.A(net13),
    .B(net51),
    .Y(_03402_));
 sky130_fd_sc_hd__nor2_1 _08987_ (.A(_03401_),
    .B(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__xnor2_1 _08988_ (.A(_03340_),
    .B(_03341_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand2_1 _08989_ (.A(net11),
    .B(net51),
    .Y(_03405_));
 sky130_fd_sc_hd__nor2_1 _08990_ (.A(_03404_),
    .B(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__xnor2_1 _08991_ (.A(_03338_),
    .B(_03339_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2_1 _08992_ (.A(net10),
    .B(net51),
    .Y(_03408_));
 sky130_fd_sc_hd__nor2_1 _08993_ (.A(_03407_),
    .B(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__xnor2_1 _08994_ (.A(_03336_),
    .B(_03337_),
    .Y(_03410_));
 sky130_fd_sc_hd__nand2_1 _08995_ (.A(net9),
    .B(net51),
    .Y(_03412_));
 sky130_fd_sc_hd__nor2_1 _08996_ (.A(_03410_),
    .B(_03412_),
    .Y(_03413_));
 sky130_fd_sc_hd__xnor2_1 _08997_ (.A(_03333_),
    .B(_03335_),
    .Y(_03414_));
 sky130_fd_sc_hd__nand2_1 _08998_ (.A(net8),
    .B(net51),
    .Y(_03415_));
 sky130_fd_sc_hd__nor2_1 _08999_ (.A(_03414_),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__xnor2_1 _09000_ (.A(_03331_),
    .B(_03332_),
    .Y(_03417_));
 sky130_fd_sc_hd__nand2_1 _09001_ (.A(net7),
    .B(net51),
    .Y(_03418_));
 sky130_fd_sc_hd__nor2_1 _09002_ (.A(_03417_),
    .B(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__xnor2_1 _09003_ (.A(_03329_),
    .B(_03330_),
    .Y(_03420_));
 sky130_fd_sc_hd__nand2_1 _09004_ (.A(net6),
    .B(net51),
    .Y(_03421_));
 sky130_fd_sc_hd__nor2_1 _09005_ (.A(_03420_),
    .B(_03421_),
    .Y(_03423_));
 sky130_fd_sc_hd__xnor2_1 _09006_ (.A(_03327_),
    .B(_03328_),
    .Y(_03424_));
 sky130_fd_sc_hd__nand2_1 _09007_ (.A(net5),
    .B(net51),
    .Y(_03425_));
 sky130_fd_sc_hd__nor2_1 _09008_ (.A(_03424_),
    .B(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__xnor2_1 _09009_ (.A(_03325_),
    .B(_03326_),
    .Y(_03427_));
 sky130_fd_sc_hd__nand2_1 _09010_ (.A(net4),
    .B(net51),
    .Y(_03428_));
 sky130_fd_sc_hd__nor2_1 _09011_ (.A(_03427_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__xnor2_1 _09012_ (.A(_03322_),
    .B(_03324_),
    .Y(_03430_));
 sky130_fd_sc_hd__nand2_1 _09013_ (.A(net3),
    .B(net51),
    .Y(_03431_));
 sky130_fd_sc_hd__nor2_1 _09014_ (.A(_03430_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__xnor2_1 _09015_ (.A(_03320_),
    .B(_03321_),
    .Y(_03434_));
 sky130_fd_sc_hd__nand2_1 _09016_ (.A(net2),
    .B(net51),
    .Y(_03435_));
 sky130_fd_sc_hd__nor2_1 _09017_ (.A(_03434_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__xnor2_1 _09018_ (.A(_03318_),
    .B(_03319_),
    .Y(_03437_));
 sky130_fd_sc_hd__nand2_1 _09019_ (.A(net32),
    .B(net51),
    .Y(_03438_));
 sky130_fd_sc_hd__nor2_1 _09020_ (.A(_03437_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__xnor2_1 _09021_ (.A(_03316_),
    .B(_03317_),
    .Y(_03440_));
 sky130_fd_sc_hd__nand2_1 _09022_ (.A(net31),
    .B(net51),
    .Y(_03441_));
 sky130_fd_sc_hd__nor2_1 _09023_ (.A(_03440_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__xnor2_1 _09024_ (.A(_03314_),
    .B(_03315_),
    .Y(_03443_));
 sky130_fd_sc_hd__nand2_1 _09025_ (.A(net30),
    .B(net51),
    .Y(_03445_));
 sky130_fd_sc_hd__nor2_1 _09026_ (.A(_03443_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__xnor2_1 _09027_ (.A(_03311_),
    .B(_03313_),
    .Y(_03447_));
 sky130_fd_sc_hd__nand2_1 _09028_ (.A(net29),
    .B(net51),
    .Y(_03448_));
 sky130_fd_sc_hd__nor2_1 _09029_ (.A(_03447_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__a21o_1 _09030_ (.A1(_01477_),
    .A2(_01618_),
    .B1(_01617_),
    .X(_03450_));
 sky130_fd_sc_hd__xor2_1 _09031_ (.A(_03447_),
    .B(_03448_),
    .X(_03451_));
 sky130_fd_sc_hd__a21o_1 _09032_ (.A1(_03450_),
    .A2(_03451_),
    .B1(_03449_),
    .X(_03452_));
 sky130_fd_sc_hd__xor2_1 _09033_ (.A(_03443_),
    .B(_03445_),
    .X(_03453_));
 sky130_fd_sc_hd__a21o_1 _09034_ (.A1(_03452_),
    .A2(_03453_),
    .B1(_03446_),
    .X(_03454_));
 sky130_fd_sc_hd__xor2_1 _09035_ (.A(_03440_),
    .B(_03441_),
    .X(_03456_));
 sky130_fd_sc_hd__a21o_1 _09036_ (.A1(_03454_),
    .A2(_03456_),
    .B1(_03442_),
    .X(_03457_));
 sky130_fd_sc_hd__xor2_1 _09037_ (.A(_03437_),
    .B(_03438_),
    .X(_03458_));
 sky130_fd_sc_hd__a21o_1 _09038_ (.A1(_03457_),
    .A2(_03458_),
    .B1(_03439_),
    .X(_03459_));
 sky130_fd_sc_hd__xor2_1 _09039_ (.A(_03434_),
    .B(_03435_),
    .X(_03460_));
 sky130_fd_sc_hd__a21o_1 _09040_ (.A1(_03459_),
    .A2(_03460_),
    .B1(_03436_),
    .X(_03461_));
 sky130_fd_sc_hd__xor2_1 _09041_ (.A(_03430_),
    .B(_03431_),
    .X(_03462_));
 sky130_fd_sc_hd__a21o_1 _09042_ (.A1(_03461_),
    .A2(_03462_),
    .B1(_03432_),
    .X(_03463_));
 sky130_fd_sc_hd__xor2_1 _09043_ (.A(_03427_),
    .B(_03428_),
    .X(_03464_));
 sky130_fd_sc_hd__a21o_1 _09044_ (.A1(_03463_),
    .A2(_03464_),
    .B1(_03429_),
    .X(_03465_));
 sky130_fd_sc_hd__xor2_1 _09045_ (.A(_03424_),
    .B(_03425_),
    .X(_03467_));
 sky130_fd_sc_hd__a21o_1 _09046_ (.A1(_03465_),
    .A2(_03467_),
    .B1(_03426_),
    .X(_03468_));
 sky130_fd_sc_hd__xor2_1 _09047_ (.A(_03420_),
    .B(_03421_),
    .X(_03469_));
 sky130_fd_sc_hd__a21o_1 _09048_ (.A1(_03468_),
    .A2(_03469_),
    .B1(_03423_),
    .X(_03470_));
 sky130_fd_sc_hd__xor2_1 _09049_ (.A(_03417_),
    .B(_03418_),
    .X(_03471_));
 sky130_fd_sc_hd__a21o_1 _09050_ (.A1(_03470_),
    .A2(_03471_),
    .B1(_03419_),
    .X(_03472_));
 sky130_fd_sc_hd__xor2_1 _09051_ (.A(_03414_),
    .B(_03415_),
    .X(_03473_));
 sky130_fd_sc_hd__a21o_1 _09052_ (.A1(_03472_),
    .A2(_03473_),
    .B1(_03416_),
    .X(_03474_));
 sky130_fd_sc_hd__xor2_1 _09053_ (.A(_03410_),
    .B(_03412_),
    .X(_03475_));
 sky130_fd_sc_hd__a21o_1 _09054_ (.A1(_03474_),
    .A2(_03475_),
    .B1(_03413_),
    .X(_03476_));
 sky130_fd_sc_hd__xor2_1 _09055_ (.A(_03407_),
    .B(_03408_),
    .X(_03478_));
 sky130_fd_sc_hd__a21o_1 _09056_ (.A1(_03476_),
    .A2(_03478_),
    .B1(_03409_),
    .X(_03479_));
 sky130_fd_sc_hd__xor2_1 _09057_ (.A(_03404_),
    .B(_03405_),
    .X(_03480_));
 sky130_fd_sc_hd__a21o_1 _09058_ (.A1(_03479_),
    .A2(_03480_),
    .B1(_03406_),
    .X(_03481_));
 sky130_fd_sc_hd__xor2_1 _09059_ (.A(_03401_),
    .B(_03402_),
    .X(_03482_));
 sky130_fd_sc_hd__a21o_1 _09060_ (.A1(_03481_),
    .A2(_03482_),
    .B1(_03403_),
    .X(_03483_));
 sky130_fd_sc_hd__xor2_1 _09061_ (.A(_03397_),
    .B(_03398_),
    .X(_03484_));
 sky130_fd_sc_hd__a21o_1 _09062_ (.A1(_03483_),
    .A2(_03484_),
    .B1(_03399_),
    .X(_03485_));
 sky130_fd_sc_hd__xor2_1 _09063_ (.A(_03394_),
    .B(_03395_),
    .X(_03486_));
 sky130_fd_sc_hd__a21o_1 _09064_ (.A1(_03485_),
    .A2(_03486_),
    .B1(_03396_),
    .X(_03487_));
 sky130_fd_sc_hd__xor2_1 _09065_ (.A(_03391_),
    .B(_03392_),
    .X(_03489_));
 sky130_fd_sc_hd__a21o_1 _09066_ (.A1(_03487_),
    .A2(_03489_),
    .B1(_03393_),
    .X(_03490_));
 sky130_fd_sc_hd__xor2_1 _09067_ (.A(_03387_),
    .B(_03388_),
    .X(_03491_));
 sky130_fd_sc_hd__a21o_1 _09068_ (.A1(_03490_),
    .A2(_03491_),
    .B1(_03390_),
    .X(_03492_));
 sky130_fd_sc_hd__xor2_1 _09069_ (.A(_03384_),
    .B(_03385_),
    .X(_03493_));
 sky130_fd_sc_hd__a21o_1 _09070_ (.A1(_03492_),
    .A2(_03493_),
    .B1(_03386_),
    .X(_03494_));
 sky130_fd_sc_hd__xor2_1 _09071_ (.A(_03381_),
    .B(_03382_),
    .X(_03495_));
 sky130_fd_sc_hd__a21o_1 _09072_ (.A1(_03494_),
    .A2(_03495_),
    .B1(_03383_),
    .X(_03496_));
 sky130_fd_sc_hd__xor2_1 _09073_ (.A(_03377_),
    .B(_03379_),
    .X(_03497_));
 sky130_fd_sc_hd__a21o_1 _09074_ (.A1(_03496_),
    .A2(_03497_),
    .B1(_03380_),
    .X(_03498_));
 sky130_fd_sc_hd__xor2_1 _09075_ (.A(_03374_),
    .B(_03375_),
    .X(_03500_));
 sky130_fd_sc_hd__a21o_1 _09076_ (.A1(_03498_),
    .A2(_03500_),
    .B1(_03376_),
    .X(_03501_));
 sky130_fd_sc_hd__xor2_1 _09077_ (.A(_03371_),
    .B(_03372_),
    .X(_03502_));
 sky130_fd_sc_hd__a21oi_1 _09078_ (.A1(_03501_),
    .A2(_03502_),
    .B1(_03373_),
    .Y(_03503_));
 sky130_fd_sc_hd__nand2_1 _09079_ (.A(net50),
    .B(net25),
    .Y(_03504_));
 sky130_fd_sc_hd__nand2_1 _09080_ (.A(_03364_),
    .B(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__or2_1 _09081_ (.A(_03364_),
    .B(_03504_),
    .X(_03506_));
 sky130_fd_sc_hd__a2bb2o_1 _09082_ (.A1_N(_03362_),
    .A2_N(_03370_),
    .B1(_03505_),
    .B2(_03506_),
    .X(_03507_));
 sky130_fd_sc_hd__a31o_1 _09083_ (.A1(net50),
    .A2(net24),
    .A3(_03368_),
    .B1(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__nand2_1 _09084_ (.A(net51),
    .B(net24),
    .Y(_03509_));
 sky130_fd_sc_hd__xor2_1 _09085_ (.A(_03508_),
    .B(_03509_),
    .X(_03511_));
 sky130_fd_sc_hd__nor2_1 _09086_ (.A(_03503_),
    .B(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__xnor2_1 _09087_ (.A(_03503_),
    .B(_03511_),
    .Y(_03513_));
 sky130_fd_sc_hd__nand2_1 _09088_ (.A(net52),
    .B(net22),
    .Y(_03514_));
 sky130_fd_sc_hd__nor2_1 _09089_ (.A(_03513_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__xnor2_1 _09090_ (.A(_03501_),
    .B(_03502_),
    .Y(_03516_));
 sky130_fd_sc_hd__nand2_1 _09091_ (.A(net52),
    .B(net21),
    .Y(_03517_));
 sky130_fd_sc_hd__nor2_1 _09092_ (.A(_03516_),
    .B(_03517_),
    .Y(_03518_));
 sky130_fd_sc_hd__xnor2_1 _09093_ (.A(_03498_),
    .B(_03500_),
    .Y(_03519_));
 sky130_fd_sc_hd__nand2_1 _09094_ (.A(net20),
    .B(net52),
    .Y(_03520_));
 sky130_fd_sc_hd__nor2_1 _09095_ (.A(_03519_),
    .B(_03520_),
    .Y(_03522_));
 sky130_fd_sc_hd__xnor2_1 _09096_ (.A(_03496_),
    .B(_03497_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand2_1 _09097_ (.A(net19),
    .B(net52),
    .Y(_03524_));
 sky130_fd_sc_hd__nor2_1 _09098_ (.A(_03523_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__xnor2_1 _09099_ (.A(_03494_),
    .B(_03495_),
    .Y(_03526_));
 sky130_fd_sc_hd__nand2_1 _09100_ (.A(net18),
    .B(net52),
    .Y(_03527_));
 sky130_fd_sc_hd__nor2_1 _09101_ (.A(_03526_),
    .B(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__xnor2_1 _09102_ (.A(_03492_),
    .B(_03493_),
    .Y(_03529_));
 sky130_fd_sc_hd__nand2_1 _09103_ (.A(net17),
    .B(net52),
    .Y(_03530_));
 sky130_fd_sc_hd__nor2_1 _09104_ (.A(_03529_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__xnor2_1 _09105_ (.A(_03490_),
    .B(_03491_),
    .Y(_03533_));
 sky130_fd_sc_hd__nand2_1 _09106_ (.A(net16),
    .B(net52),
    .Y(_03534_));
 sky130_fd_sc_hd__nor2_1 _09107_ (.A(_03533_),
    .B(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__xnor2_1 _09108_ (.A(_03487_),
    .B(_03489_),
    .Y(_03536_));
 sky130_fd_sc_hd__nand2_1 _09109_ (.A(net15),
    .B(net52),
    .Y(_03537_));
 sky130_fd_sc_hd__nor2_1 _09110_ (.A(_03536_),
    .B(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__xnor2_1 _09111_ (.A(_03485_),
    .B(_03486_),
    .Y(_03539_));
 sky130_fd_sc_hd__nand2_1 _09112_ (.A(net14),
    .B(net52),
    .Y(_03540_));
 sky130_fd_sc_hd__nor2_1 _09113_ (.A(_03539_),
    .B(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__xnor2_1 _09114_ (.A(_03483_),
    .B(_03484_),
    .Y(_03542_));
 sky130_fd_sc_hd__nand2_1 _09115_ (.A(net13),
    .B(net52),
    .Y(_03544_));
 sky130_fd_sc_hd__nor2_1 _09116_ (.A(_03542_),
    .B(_03544_),
    .Y(_03545_));
 sky130_fd_sc_hd__xnor2_1 _09117_ (.A(_03481_),
    .B(_03482_),
    .Y(_03546_));
 sky130_fd_sc_hd__nand2_1 _09118_ (.A(net11),
    .B(net52),
    .Y(_03547_));
 sky130_fd_sc_hd__nor2_1 _09119_ (.A(_03546_),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__xnor2_1 _09120_ (.A(_03479_),
    .B(_03480_),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_1 _09121_ (.A(net10),
    .B(net52),
    .Y(_03550_));
 sky130_fd_sc_hd__nor2_1 _09122_ (.A(_03549_),
    .B(_03550_),
    .Y(_03551_));
 sky130_fd_sc_hd__xnor2_1 _09123_ (.A(_03476_),
    .B(_03478_),
    .Y(_03552_));
 sky130_fd_sc_hd__nand2_1 _09124_ (.A(net9),
    .B(net52),
    .Y(_03553_));
 sky130_fd_sc_hd__nor2_1 _09125_ (.A(_03552_),
    .B(_03553_),
    .Y(_03555_));
 sky130_fd_sc_hd__xnor2_1 _09126_ (.A(_03474_),
    .B(_03475_),
    .Y(_03556_));
 sky130_fd_sc_hd__nand2_1 _09127_ (.A(net8),
    .B(net52),
    .Y(_03557_));
 sky130_fd_sc_hd__nor2_1 _09128_ (.A(_03556_),
    .B(_03557_),
    .Y(_03558_));
 sky130_fd_sc_hd__xnor2_1 _09129_ (.A(_03472_),
    .B(_03473_),
    .Y(_03559_));
 sky130_fd_sc_hd__nand2_1 _09130_ (.A(net7),
    .B(net52),
    .Y(_03560_));
 sky130_fd_sc_hd__nor2_1 _09131_ (.A(_03559_),
    .B(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__xnor2_1 _09132_ (.A(_03470_),
    .B(_03471_),
    .Y(_03562_));
 sky130_fd_sc_hd__nand2_1 _09133_ (.A(net6),
    .B(net52),
    .Y(_03563_));
 sky130_fd_sc_hd__nor2_1 _09134_ (.A(_03562_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__xnor2_1 _09135_ (.A(_03468_),
    .B(_03469_),
    .Y(_03566_));
 sky130_fd_sc_hd__nand2_1 _09136_ (.A(net5),
    .B(net52),
    .Y(_03567_));
 sky130_fd_sc_hd__nor2_1 _09137_ (.A(_03566_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__xnor2_1 _09138_ (.A(_03465_),
    .B(_03467_),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _09139_ (.A(net4),
    .B(net52),
    .Y(_03570_));
 sky130_fd_sc_hd__nor2_1 _09140_ (.A(_03569_),
    .B(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__xnor2_1 _09141_ (.A(_03463_),
    .B(_03464_),
    .Y(_03572_));
 sky130_fd_sc_hd__nand2_1 _09142_ (.A(net3),
    .B(net52),
    .Y(_03573_));
 sky130_fd_sc_hd__nor2_1 _09143_ (.A(_03572_),
    .B(_03573_),
    .Y(_03574_));
 sky130_fd_sc_hd__xnor2_1 _09144_ (.A(_03461_),
    .B(_03462_),
    .Y(_03575_));
 sky130_fd_sc_hd__nand2_1 _09145_ (.A(net2),
    .B(net52),
    .Y(_03577_));
 sky130_fd_sc_hd__nor2_1 _09146_ (.A(_03575_),
    .B(_03577_),
    .Y(_03578_));
 sky130_fd_sc_hd__xnor2_1 _09147_ (.A(_03459_),
    .B(_03460_),
    .Y(_03579_));
 sky130_fd_sc_hd__nand2_1 _09148_ (.A(net32),
    .B(net52),
    .Y(_03580_));
 sky130_fd_sc_hd__nor2_1 _09149_ (.A(_03579_),
    .B(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__xnor2_1 _09150_ (.A(_03457_),
    .B(_03458_),
    .Y(_03582_));
 sky130_fd_sc_hd__nand2_1 _09151_ (.A(net31),
    .B(net52),
    .Y(_03583_));
 sky130_fd_sc_hd__nor2_1 _09152_ (.A(_03582_),
    .B(_03583_),
    .Y(_03584_));
 sky130_fd_sc_hd__xnor2_1 _09153_ (.A(_03454_),
    .B(_03456_),
    .Y(_03585_));
 sky130_fd_sc_hd__nand2_1 _09154_ (.A(net30),
    .B(net52),
    .Y(_03586_));
 sky130_fd_sc_hd__nor2_1 _09155_ (.A(_03585_),
    .B(_03586_),
    .Y(_03588_));
 sky130_fd_sc_hd__xnor2_1 _09156_ (.A(_03452_),
    .B(_03453_),
    .Y(_03589_));
 sky130_fd_sc_hd__nand2_1 _09157_ (.A(net29),
    .B(net52),
    .Y(_03590_));
 sky130_fd_sc_hd__nor2_1 _09158_ (.A(_03589_),
    .B(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__xnor2_1 _09159_ (.A(_03450_),
    .B(_03451_),
    .Y(_03592_));
 sky130_fd_sc_hd__nand2_1 _09160_ (.A(net28),
    .B(net52),
    .Y(_03593_));
 sky130_fd_sc_hd__nor2_1 _09161_ (.A(_03592_),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__a21o_1 _09162_ (.A1(_01474_),
    .A2(_01622_),
    .B1(_01621_),
    .X(_03595_));
 sky130_fd_sc_hd__xor2_1 _09163_ (.A(_03592_),
    .B(_03593_),
    .X(_03596_));
 sky130_fd_sc_hd__a21o_1 _09164_ (.A1(_03595_),
    .A2(_03596_),
    .B1(_03594_),
    .X(_03597_));
 sky130_fd_sc_hd__xor2_1 _09165_ (.A(_03589_),
    .B(_03590_),
    .X(_03599_));
 sky130_fd_sc_hd__a21o_1 _09166_ (.A1(_03597_),
    .A2(_03599_),
    .B1(_03591_),
    .X(_03600_));
 sky130_fd_sc_hd__xor2_1 _09167_ (.A(_03585_),
    .B(_03586_),
    .X(_03601_));
 sky130_fd_sc_hd__a21o_1 _09168_ (.A1(_03600_),
    .A2(_03601_),
    .B1(_03588_),
    .X(_03602_));
 sky130_fd_sc_hd__xor2_1 _09169_ (.A(_03582_),
    .B(_03583_),
    .X(_03603_));
 sky130_fd_sc_hd__a21o_1 _09170_ (.A1(_03602_),
    .A2(_03603_),
    .B1(_03584_),
    .X(_03604_));
 sky130_fd_sc_hd__xor2_1 _09171_ (.A(_03579_),
    .B(_03580_),
    .X(_03605_));
 sky130_fd_sc_hd__a21o_1 _09172_ (.A1(_03604_),
    .A2(_03605_),
    .B1(_03581_),
    .X(_03606_));
 sky130_fd_sc_hd__xor2_1 _09173_ (.A(_03575_),
    .B(_03577_),
    .X(_03607_));
 sky130_fd_sc_hd__a21o_1 _09174_ (.A1(_03606_),
    .A2(_03607_),
    .B1(_03578_),
    .X(_03608_));
 sky130_fd_sc_hd__xor2_1 _09175_ (.A(_03572_),
    .B(_03573_),
    .X(_03610_));
 sky130_fd_sc_hd__a21o_1 _09176_ (.A1(_03608_),
    .A2(_03610_),
    .B1(_03574_),
    .X(_03611_));
 sky130_fd_sc_hd__xor2_1 _09177_ (.A(_03569_),
    .B(_03570_),
    .X(_03612_));
 sky130_fd_sc_hd__a21o_1 _09178_ (.A1(_03611_),
    .A2(_03612_),
    .B1(_03571_),
    .X(_03613_));
 sky130_fd_sc_hd__xor2_1 _09179_ (.A(_03566_),
    .B(_03567_),
    .X(_03614_));
 sky130_fd_sc_hd__a21o_1 _09180_ (.A1(_03613_),
    .A2(_03614_),
    .B1(_03568_),
    .X(_03615_));
 sky130_fd_sc_hd__xor2_1 _09181_ (.A(_03562_),
    .B(_03563_),
    .X(_03616_));
 sky130_fd_sc_hd__a21o_1 _09182_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_03564_),
    .X(_03617_));
 sky130_fd_sc_hd__xor2_1 _09183_ (.A(_03559_),
    .B(_03560_),
    .X(_03618_));
 sky130_fd_sc_hd__a21o_1 _09184_ (.A1(_03617_),
    .A2(_03618_),
    .B1(_03561_),
    .X(_03619_));
 sky130_fd_sc_hd__xor2_1 _09185_ (.A(_03556_),
    .B(_03557_),
    .X(_03621_));
 sky130_fd_sc_hd__a21o_1 _09186_ (.A1(_03619_),
    .A2(_03621_),
    .B1(_03558_),
    .X(_03622_));
 sky130_fd_sc_hd__xor2_1 _09187_ (.A(_03552_),
    .B(_03553_),
    .X(_03623_));
 sky130_fd_sc_hd__a21o_1 _09188_ (.A1(_03622_),
    .A2(_03623_),
    .B1(_03555_),
    .X(_03624_));
 sky130_fd_sc_hd__xor2_1 _09189_ (.A(_03549_),
    .B(_03550_),
    .X(_03625_));
 sky130_fd_sc_hd__a21o_1 _09190_ (.A1(_03624_),
    .A2(_03625_),
    .B1(_03551_),
    .X(_03626_));
 sky130_fd_sc_hd__xor2_1 _09191_ (.A(_03546_),
    .B(_03547_),
    .X(_03627_));
 sky130_fd_sc_hd__a21o_1 _09192_ (.A1(_03626_),
    .A2(_03627_),
    .B1(_03548_),
    .X(_03628_));
 sky130_fd_sc_hd__xor2_1 _09193_ (.A(_03542_),
    .B(_03544_),
    .X(_03629_));
 sky130_fd_sc_hd__a21o_1 _09194_ (.A1(_03628_),
    .A2(_03629_),
    .B1(_03545_),
    .X(_03630_));
 sky130_fd_sc_hd__xor2_1 _09195_ (.A(_03539_),
    .B(_03540_),
    .X(_03632_));
 sky130_fd_sc_hd__a21o_1 _09196_ (.A1(_03630_),
    .A2(_03632_),
    .B1(_03541_),
    .X(_03633_));
 sky130_fd_sc_hd__xor2_1 _09197_ (.A(_03536_),
    .B(_03537_),
    .X(_03634_));
 sky130_fd_sc_hd__a21o_1 _09198_ (.A1(_03633_),
    .A2(_03634_),
    .B1(_03538_),
    .X(_03635_));
 sky130_fd_sc_hd__xor2_1 _09199_ (.A(_03533_),
    .B(_03534_),
    .X(_03636_));
 sky130_fd_sc_hd__a21o_1 _09200_ (.A1(_03635_),
    .A2(_03636_),
    .B1(_03535_),
    .X(_03637_));
 sky130_fd_sc_hd__xor2_1 _09201_ (.A(_03529_),
    .B(_03530_),
    .X(_03638_));
 sky130_fd_sc_hd__a21o_1 _09202_ (.A1(_03637_),
    .A2(_03638_),
    .B1(_03531_),
    .X(_03639_));
 sky130_fd_sc_hd__xor2_1 _09203_ (.A(_03526_),
    .B(_03527_),
    .X(_03640_));
 sky130_fd_sc_hd__a21o_1 _09204_ (.A1(_03639_),
    .A2(_03640_),
    .B1(_03528_),
    .X(_03641_));
 sky130_fd_sc_hd__xor2_1 _09205_ (.A(_03523_),
    .B(_03524_),
    .X(_03643_));
 sky130_fd_sc_hd__a21o_1 _09206_ (.A1(_03641_),
    .A2(_03643_),
    .B1(_03525_),
    .X(_03644_));
 sky130_fd_sc_hd__xor2_1 _09207_ (.A(_03519_),
    .B(_03520_),
    .X(_03645_));
 sky130_fd_sc_hd__a21o_1 _09208_ (.A1(_03644_),
    .A2(_03645_),
    .B1(_03522_),
    .X(_03646_));
 sky130_fd_sc_hd__xor2_1 _09209_ (.A(_03516_),
    .B(_03517_),
    .X(_03647_));
 sky130_fd_sc_hd__a21o_1 _09210_ (.A1(_03646_),
    .A2(_03647_),
    .B1(_03518_),
    .X(_03648_));
 sky130_fd_sc_hd__xor2_1 _09211_ (.A(_03513_),
    .B(_03514_),
    .X(_03649_));
 sky130_fd_sc_hd__a21oi_1 _09212_ (.A1(_03648_),
    .A2(_03649_),
    .B1(_03515_),
    .Y(_03650_));
 sky130_fd_sc_hd__nand2_1 _09213_ (.A(net51),
    .B(net25),
    .Y(_03651_));
 sky130_fd_sc_hd__and3_1 _09214_ (.A(_03364_),
    .B(_03504_),
    .C(_03651_),
    .X(_03652_));
 sky130_fd_sc_hd__and3_1 _09215_ (.A(net51),
    .B(net25),
    .C(_03505_),
    .X(_03654_));
 sky130_fd_sc_hd__nor2_1 _09216_ (.A(_03652_),
    .B(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__a311o_1 _09217_ (.A1(net51),
    .A2(net24),
    .A3(_03508_),
    .B1(_03512_),
    .C1(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__nand2_1 _09218_ (.A(net52),
    .B(net24),
    .Y(_03657_));
 sky130_fd_sc_hd__xor2_1 _09219_ (.A(_03656_),
    .B(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__xnor2_1 _09220_ (.A(_03650_),
    .B(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__nand2_1 _09221_ (.A(net53),
    .B(net22),
    .Y(_03660_));
 sky130_fd_sc_hd__nor2_1 _09222_ (.A(_03659_),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__xnor2_1 _09223_ (.A(_03648_),
    .B(_03649_),
    .Y(_03662_));
 sky130_fd_sc_hd__nand2_1 _09224_ (.A(net21),
    .B(net53),
    .Y(_03663_));
 sky130_fd_sc_hd__nor2_1 _09225_ (.A(_03662_),
    .B(_03663_),
    .Y(_03665_));
 sky130_fd_sc_hd__xnor2_1 _09226_ (.A(_03646_),
    .B(_03647_),
    .Y(_03666_));
 sky130_fd_sc_hd__nand2_1 _09227_ (.A(net20),
    .B(net53),
    .Y(_03667_));
 sky130_fd_sc_hd__nor2_1 _09228_ (.A(_03666_),
    .B(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__xnor2_1 _09229_ (.A(_03644_),
    .B(_03645_),
    .Y(_03669_));
 sky130_fd_sc_hd__nand2_1 _09230_ (.A(net19),
    .B(net53),
    .Y(_03670_));
 sky130_fd_sc_hd__nor2_1 _09231_ (.A(_03669_),
    .B(_03670_),
    .Y(_03671_));
 sky130_fd_sc_hd__xnor2_1 _09232_ (.A(_03641_),
    .B(_03643_),
    .Y(_03672_));
 sky130_fd_sc_hd__nand2_1 _09233_ (.A(net18),
    .B(net53),
    .Y(_03673_));
 sky130_fd_sc_hd__nor2_1 _09234_ (.A(_03672_),
    .B(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__xnor2_1 _09235_ (.A(_03639_),
    .B(_03640_),
    .Y(_03676_));
 sky130_fd_sc_hd__nand2_1 _09236_ (.A(net17),
    .B(net53),
    .Y(_03677_));
 sky130_fd_sc_hd__nor2_1 _09237_ (.A(_03676_),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__xnor2_1 _09238_ (.A(_03637_),
    .B(_03638_),
    .Y(_03679_));
 sky130_fd_sc_hd__nand2_1 _09239_ (.A(net16),
    .B(net53),
    .Y(_03680_));
 sky130_fd_sc_hd__nor2_1 _09240_ (.A(_03679_),
    .B(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__xnor2_1 _09241_ (.A(_03635_),
    .B(_03636_),
    .Y(_03682_));
 sky130_fd_sc_hd__nand2_1 _09242_ (.A(net15),
    .B(net53),
    .Y(_03683_));
 sky130_fd_sc_hd__nor2_1 _09243_ (.A(_03682_),
    .B(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__xnor2_1 _09244_ (.A(_03633_),
    .B(_03634_),
    .Y(_03685_));
 sky130_fd_sc_hd__nand2_1 _09245_ (.A(net14),
    .B(net53),
    .Y(_03687_));
 sky130_fd_sc_hd__nor2_1 _09246_ (.A(_03685_),
    .B(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__xnor2_1 _09247_ (.A(_03630_),
    .B(_03632_),
    .Y(_03689_));
 sky130_fd_sc_hd__nand2_1 _09248_ (.A(net13),
    .B(net53),
    .Y(_03690_));
 sky130_fd_sc_hd__nor2_1 _09249_ (.A(_03689_),
    .B(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__xnor2_1 _09250_ (.A(_03628_),
    .B(_03629_),
    .Y(_03692_));
 sky130_fd_sc_hd__nand2_1 _09251_ (.A(net11),
    .B(net53),
    .Y(_03693_));
 sky130_fd_sc_hd__nor2_1 _09252_ (.A(_03692_),
    .B(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__xnor2_1 _09253_ (.A(_03626_),
    .B(_03627_),
    .Y(_03695_));
 sky130_fd_sc_hd__nand2_1 _09254_ (.A(net10),
    .B(net53),
    .Y(_03696_));
 sky130_fd_sc_hd__nor2_1 _09255_ (.A(_03695_),
    .B(_03696_),
    .Y(_03698_));
 sky130_fd_sc_hd__xnor2_1 _09256_ (.A(_03624_),
    .B(_03625_),
    .Y(_03699_));
 sky130_fd_sc_hd__nand2_1 _09257_ (.A(net9),
    .B(net53),
    .Y(_03700_));
 sky130_fd_sc_hd__nor2_1 _09258_ (.A(_03699_),
    .B(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__xnor2_1 _09259_ (.A(_03622_),
    .B(_03623_),
    .Y(_03702_));
 sky130_fd_sc_hd__nand2_1 _09260_ (.A(net8),
    .B(net53),
    .Y(_03703_));
 sky130_fd_sc_hd__nor2_1 _09261_ (.A(_03702_),
    .B(_03703_),
    .Y(_03704_));
 sky130_fd_sc_hd__xnor2_1 _09262_ (.A(_03619_),
    .B(_03621_),
    .Y(_03705_));
 sky130_fd_sc_hd__nand2_1 _09263_ (.A(net7),
    .B(net53),
    .Y(_03706_));
 sky130_fd_sc_hd__nor2_1 _09264_ (.A(_03705_),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__xnor2_1 _09265_ (.A(_03617_),
    .B(_03618_),
    .Y(_03709_));
 sky130_fd_sc_hd__nand2_1 _09266_ (.A(net6),
    .B(net53),
    .Y(_03710_));
 sky130_fd_sc_hd__nor2_1 _09267_ (.A(_03709_),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__xnor2_1 _09268_ (.A(_03615_),
    .B(_03616_),
    .Y(_03712_));
 sky130_fd_sc_hd__nand2_1 _09269_ (.A(net5),
    .B(net53),
    .Y(_03713_));
 sky130_fd_sc_hd__nor2_1 _09270_ (.A(_03712_),
    .B(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__xnor2_1 _09271_ (.A(_03613_),
    .B(_03614_),
    .Y(_03715_));
 sky130_fd_sc_hd__nand2_1 _09272_ (.A(net4),
    .B(net53),
    .Y(_03716_));
 sky130_fd_sc_hd__nor2_1 _09273_ (.A(_03715_),
    .B(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__xnor2_1 _09274_ (.A(_03611_),
    .B(_03612_),
    .Y(_03718_));
 sky130_fd_sc_hd__nand2_1 _09275_ (.A(net3),
    .B(net53),
    .Y(_03720_));
 sky130_fd_sc_hd__nor2_1 _09276_ (.A(_03718_),
    .B(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__xnor2_1 _09277_ (.A(_03608_),
    .B(_03610_),
    .Y(_03722_));
 sky130_fd_sc_hd__nand2_1 _09278_ (.A(net2),
    .B(net53),
    .Y(_03723_));
 sky130_fd_sc_hd__nor2_1 _09279_ (.A(_03722_),
    .B(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__xnor2_1 _09280_ (.A(_03606_),
    .B(_03607_),
    .Y(_03725_));
 sky130_fd_sc_hd__nand2_1 _09281_ (.A(net32),
    .B(net53),
    .Y(_03726_));
 sky130_fd_sc_hd__nor2_1 _09282_ (.A(_03725_),
    .B(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__xnor2_1 _09283_ (.A(_03604_),
    .B(_03605_),
    .Y(_03728_));
 sky130_fd_sc_hd__nand2_1 _09284_ (.A(net31),
    .B(net53),
    .Y(_03729_));
 sky130_fd_sc_hd__nor2_1 _09285_ (.A(_03728_),
    .B(_03729_),
    .Y(_03731_));
 sky130_fd_sc_hd__xnor2_1 _09286_ (.A(_03602_),
    .B(_03603_),
    .Y(_03732_));
 sky130_fd_sc_hd__nand2_1 _09287_ (.A(net30),
    .B(net53),
    .Y(_03733_));
 sky130_fd_sc_hd__nor2_1 _09288_ (.A(_03732_),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__xnor2_1 _09289_ (.A(_03600_),
    .B(_03601_),
    .Y(_03735_));
 sky130_fd_sc_hd__nand2_1 _09290_ (.A(net29),
    .B(net53),
    .Y(_03736_));
 sky130_fd_sc_hd__nor2_1 _09291_ (.A(_03735_),
    .B(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__xnor2_1 _09292_ (.A(_03597_),
    .B(_03599_),
    .Y(_03738_));
 sky130_fd_sc_hd__nand2_1 _09293_ (.A(net28),
    .B(net53),
    .Y(_03739_));
 sky130_fd_sc_hd__nor2_1 _09294_ (.A(_03738_),
    .B(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__xnor2_1 _09295_ (.A(_03595_),
    .B(_03596_),
    .Y(_03742_));
 sky130_fd_sc_hd__nand2_1 _09296_ (.A(net27),
    .B(net53),
    .Y(_03743_));
 sky130_fd_sc_hd__nor2_1 _09297_ (.A(_03742_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__a21o_1 _09298_ (.A1(_01472_),
    .A2(_01625_),
    .B1(_01624_),
    .X(_03745_));
 sky130_fd_sc_hd__xor2_1 _09299_ (.A(_03742_),
    .B(_03743_),
    .X(_03746_));
 sky130_fd_sc_hd__a21o_1 _09300_ (.A1(_03745_),
    .A2(_03746_),
    .B1(_03744_),
    .X(_03747_));
 sky130_fd_sc_hd__xor2_1 _09301_ (.A(_03738_),
    .B(_03739_),
    .X(_03748_));
 sky130_fd_sc_hd__a21o_1 _09302_ (.A1(_03747_),
    .A2(_03748_),
    .B1(_03740_),
    .X(_03749_));
 sky130_fd_sc_hd__xor2_1 _09303_ (.A(_03735_),
    .B(_03736_),
    .X(_03750_));
 sky130_fd_sc_hd__a21o_1 _09304_ (.A1(_03749_),
    .A2(_03750_),
    .B1(_03737_),
    .X(_03751_));
 sky130_fd_sc_hd__xor2_1 _09305_ (.A(_03732_),
    .B(_03733_),
    .X(_03753_));
 sky130_fd_sc_hd__a21o_1 _09306_ (.A1(_03751_),
    .A2(_03753_),
    .B1(_03734_),
    .X(_03754_));
 sky130_fd_sc_hd__xor2_1 _09307_ (.A(_03728_),
    .B(_03729_),
    .X(_03755_));
 sky130_fd_sc_hd__a21o_1 _09308_ (.A1(_03754_),
    .A2(_03755_),
    .B1(_03731_),
    .X(_03756_));
 sky130_fd_sc_hd__xor2_1 _09309_ (.A(_03725_),
    .B(_03726_),
    .X(_03757_));
 sky130_fd_sc_hd__a21o_1 _09310_ (.A1(_03756_),
    .A2(_03757_),
    .B1(_03727_),
    .X(_03758_));
 sky130_fd_sc_hd__xor2_1 _09311_ (.A(_03722_),
    .B(_03723_),
    .X(_03759_));
 sky130_fd_sc_hd__a21o_1 _09312_ (.A1(_03758_),
    .A2(_03759_),
    .B1(_03724_),
    .X(_03760_));
 sky130_fd_sc_hd__xor2_1 _09313_ (.A(_03718_),
    .B(_03720_),
    .X(_03761_));
 sky130_fd_sc_hd__a21o_1 _09314_ (.A1(_03760_),
    .A2(_03761_),
    .B1(_03721_),
    .X(_03762_));
 sky130_fd_sc_hd__xor2_1 _09315_ (.A(_03715_),
    .B(_03716_),
    .X(_03764_));
 sky130_fd_sc_hd__a21o_1 _09316_ (.A1(_03762_),
    .A2(_03764_),
    .B1(_03717_),
    .X(_03765_));
 sky130_fd_sc_hd__xor2_1 _09317_ (.A(_03712_),
    .B(_03713_),
    .X(_03766_));
 sky130_fd_sc_hd__a21o_1 _09318_ (.A1(_03765_),
    .A2(_03766_),
    .B1(_03714_),
    .X(_03767_));
 sky130_fd_sc_hd__xor2_1 _09319_ (.A(_03709_),
    .B(_03710_),
    .X(_03768_));
 sky130_fd_sc_hd__a21o_1 _09320_ (.A1(_03767_),
    .A2(_03768_),
    .B1(_03711_),
    .X(_03769_));
 sky130_fd_sc_hd__xor2_1 _09321_ (.A(_03705_),
    .B(_03706_),
    .X(_03770_));
 sky130_fd_sc_hd__a21o_1 _09322_ (.A1(_03769_),
    .A2(_03770_),
    .B1(_03707_),
    .X(_03771_));
 sky130_fd_sc_hd__xor2_1 _09323_ (.A(_03702_),
    .B(_03703_),
    .X(_03772_));
 sky130_fd_sc_hd__a21o_1 _09324_ (.A1(_03771_),
    .A2(_03772_),
    .B1(_03704_),
    .X(_03773_));
 sky130_fd_sc_hd__xor2_1 _09325_ (.A(_03699_),
    .B(_03700_),
    .X(_03775_));
 sky130_fd_sc_hd__a21o_1 _09326_ (.A1(_03773_),
    .A2(_03775_),
    .B1(_03701_),
    .X(_03776_));
 sky130_fd_sc_hd__xor2_1 _09327_ (.A(_03695_),
    .B(_03696_),
    .X(_03777_));
 sky130_fd_sc_hd__a21o_1 _09328_ (.A1(_03776_),
    .A2(_03777_),
    .B1(_03698_),
    .X(_03778_));
 sky130_fd_sc_hd__xor2_1 _09329_ (.A(_03692_),
    .B(_03693_),
    .X(_03779_));
 sky130_fd_sc_hd__a21o_1 _09330_ (.A1(_03778_),
    .A2(_03779_),
    .B1(_03694_),
    .X(_03780_));
 sky130_fd_sc_hd__xor2_1 _09331_ (.A(_03689_),
    .B(_03690_),
    .X(_03781_));
 sky130_fd_sc_hd__a21o_1 _09332_ (.A1(_03780_),
    .A2(_03781_),
    .B1(_03691_),
    .X(_03782_));
 sky130_fd_sc_hd__xor2_1 _09333_ (.A(_03685_),
    .B(_03687_),
    .X(_03783_));
 sky130_fd_sc_hd__a21o_1 _09334_ (.A1(_03782_),
    .A2(_03783_),
    .B1(_03688_),
    .X(_03784_));
 sky130_fd_sc_hd__xor2_1 _09335_ (.A(_03682_),
    .B(_03683_),
    .X(_03786_));
 sky130_fd_sc_hd__a21o_1 _09336_ (.A1(_03784_),
    .A2(_03786_),
    .B1(_03684_),
    .X(_03787_));
 sky130_fd_sc_hd__xor2_1 _09337_ (.A(_03679_),
    .B(_03680_),
    .X(_03788_));
 sky130_fd_sc_hd__a21o_1 _09338_ (.A1(_03787_),
    .A2(_03788_),
    .B1(_03681_),
    .X(_03789_));
 sky130_fd_sc_hd__xor2_1 _09339_ (.A(_03676_),
    .B(_03677_),
    .X(_03790_));
 sky130_fd_sc_hd__a21o_1 _09340_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03678_),
    .X(_03791_));
 sky130_fd_sc_hd__xor2_1 _09341_ (.A(_03672_),
    .B(_03673_),
    .X(_03792_));
 sky130_fd_sc_hd__a21o_1 _09342_ (.A1(_03791_),
    .A2(_03792_),
    .B1(_03674_),
    .X(_03793_));
 sky130_fd_sc_hd__xor2_1 _09343_ (.A(_03669_),
    .B(_03670_),
    .X(_03794_));
 sky130_fd_sc_hd__a21o_1 _09344_ (.A1(_03793_),
    .A2(_03794_),
    .B1(_03671_),
    .X(_03795_));
 sky130_fd_sc_hd__xor2_1 _09345_ (.A(_03666_),
    .B(_03667_),
    .X(_03797_));
 sky130_fd_sc_hd__a21o_1 _09346_ (.A1(_03795_),
    .A2(_03797_),
    .B1(_03668_),
    .X(_03798_));
 sky130_fd_sc_hd__xor2_1 _09347_ (.A(_03662_),
    .B(_03663_),
    .X(_03799_));
 sky130_fd_sc_hd__a21o_1 _09348_ (.A1(_03798_),
    .A2(_03799_),
    .B1(_03665_),
    .X(_03800_));
 sky130_fd_sc_hd__xor2_1 _09349_ (.A(_03659_),
    .B(_03660_),
    .X(_03801_));
 sky130_fd_sc_hd__a21oi_1 _09350_ (.A1(_03800_),
    .A2(_03801_),
    .B1(_03661_),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_1 _09351_ (.A(net52),
    .B(net25),
    .Y(_03803_));
 sky130_fd_sc_hd__nand2_1 _09352_ (.A(_03652_),
    .B(_03803_),
    .Y(_03804_));
 sky130_fd_sc_hd__or2_1 _09353_ (.A(_03652_),
    .B(_03803_),
    .X(_03805_));
 sky130_fd_sc_hd__a2bb2o_1 _09354_ (.A1_N(_03650_),
    .A2_N(_03658_),
    .B1(_03804_),
    .B2(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__a31o_1 _09355_ (.A1(net52),
    .A2(net24),
    .A3(_03656_),
    .B1(_03806_),
    .X(_03808_));
 sky130_fd_sc_hd__nand2_1 _09356_ (.A(net53),
    .B(net24),
    .Y(_03809_));
 sky130_fd_sc_hd__and3_1 _09357_ (.A(net53),
    .B(net24),
    .C(_03808_),
    .X(_03810_));
 sky130_fd_sc_hd__xor2_1 _09358_ (.A(_03808_),
    .B(_03809_),
    .X(_03811_));
 sky130_fd_sc_hd__nor2_1 _09359_ (.A(_03802_),
    .B(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hd__xnor2_1 _09360_ (.A(_03802_),
    .B(_03811_),
    .Y(_03813_));
 sky130_fd_sc_hd__nand2_1 _09361_ (.A(net22),
    .B(net54),
    .Y(_03814_));
 sky130_fd_sc_hd__nor2_1 _09362_ (.A(_03813_),
    .B(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__xnor2_1 _09363_ (.A(_03800_),
    .B(_03801_),
    .Y(_03816_));
 sky130_fd_sc_hd__nand2_1 _09364_ (.A(net21),
    .B(net54),
    .Y(_03817_));
 sky130_fd_sc_hd__nor2_1 _09365_ (.A(_03816_),
    .B(_03817_),
    .Y(_03819_));
 sky130_fd_sc_hd__xnor2_1 _09366_ (.A(_03798_),
    .B(_03799_),
    .Y(_03820_));
 sky130_fd_sc_hd__nand2_1 _09367_ (.A(net20),
    .B(net54),
    .Y(_03821_));
 sky130_fd_sc_hd__nor2_1 _09368_ (.A(_03820_),
    .B(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__xnor2_1 _09369_ (.A(_03795_),
    .B(_03797_),
    .Y(_03823_));
 sky130_fd_sc_hd__nand2_1 _09370_ (.A(net19),
    .B(net54),
    .Y(_03824_));
 sky130_fd_sc_hd__nor2_1 _09371_ (.A(_03823_),
    .B(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__xnor2_1 _09372_ (.A(_03793_),
    .B(_03794_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand2_1 _09373_ (.A(net18),
    .B(net54),
    .Y(_03827_));
 sky130_fd_sc_hd__nor2_1 _09374_ (.A(_03826_),
    .B(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__xnor2_1 _09375_ (.A(_03791_),
    .B(_03792_),
    .Y(_03830_));
 sky130_fd_sc_hd__nand2_1 _09376_ (.A(net17),
    .B(net54),
    .Y(_03831_));
 sky130_fd_sc_hd__nor2_1 _09377_ (.A(_03830_),
    .B(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__xnor2_1 _09378_ (.A(_03789_),
    .B(_03790_),
    .Y(_03833_));
 sky130_fd_sc_hd__nand2_1 _09379_ (.A(net16),
    .B(net54),
    .Y(_03834_));
 sky130_fd_sc_hd__nor2_1 _09380_ (.A(_03833_),
    .B(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__xnor2_1 _09381_ (.A(_03787_),
    .B(_03788_),
    .Y(_03836_));
 sky130_fd_sc_hd__nand2_1 _09382_ (.A(net15),
    .B(net54),
    .Y(_03837_));
 sky130_fd_sc_hd__nor2_1 _09383_ (.A(_03836_),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__xnor2_1 _09384_ (.A(_03784_),
    .B(_03786_),
    .Y(_03839_));
 sky130_fd_sc_hd__nand2_1 _09385_ (.A(net14),
    .B(net54),
    .Y(_03841_));
 sky130_fd_sc_hd__nor2_1 _09386_ (.A(_03839_),
    .B(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__xnor2_1 _09387_ (.A(_03782_),
    .B(_03783_),
    .Y(_03843_));
 sky130_fd_sc_hd__nand2_1 _09388_ (.A(net13),
    .B(net54),
    .Y(_03844_));
 sky130_fd_sc_hd__nor2_1 _09389_ (.A(_03843_),
    .B(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__xnor2_1 _09390_ (.A(_03780_),
    .B(_03781_),
    .Y(_03846_));
 sky130_fd_sc_hd__nand2_1 _09391_ (.A(net11),
    .B(net54),
    .Y(_03847_));
 sky130_fd_sc_hd__nor2_1 _09392_ (.A(_03846_),
    .B(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__xnor2_1 _09393_ (.A(_03778_),
    .B(_03779_),
    .Y(_03849_));
 sky130_fd_sc_hd__nand2_1 _09394_ (.A(net10),
    .B(net54),
    .Y(_03850_));
 sky130_fd_sc_hd__nor2_1 _09395_ (.A(_03849_),
    .B(_03850_),
    .Y(_03852_));
 sky130_fd_sc_hd__xnor2_1 _09396_ (.A(_03776_),
    .B(_03777_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2_1 _09397_ (.A(net9),
    .B(net54),
    .Y(_03854_));
 sky130_fd_sc_hd__nor2_1 _09398_ (.A(_03853_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__xnor2_1 _09399_ (.A(_03773_),
    .B(_03775_),
    .Y(_03856_));
 sky130_fd_sc_hd__nand2_1 _09400_ (.A(net8),
    .B(net54),
    .Y(_03857_));
 sky130_fd_sc_hd__nor2_1 _09401_ (.A(_03856_),
    .B(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__xnor2_1 _09402_ (.A(_03771_),
    .B(_03772_),
    .Y(_03859_));
 sky130_fd_sc_hd__nand2_1 _09403_ (.A(net7),
    .B(net54),
    .Y(_03860_));
 sky130_fd_sc_hd__nor2_1 _09404_ (.A(_03859_),
    .B(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__xnor2_1 _09405_ (.A(_03769_),
    .B(_03770_),
    .Y(_03863_));
 sky130_fd_sc_hd__nand2_1 _09406_ (.A(net6),
    .B(net54),
    .Y(_03864_));
 sky130_fd_sc_hd__nor2_1 _09407_ (.A(_03863_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__xnor2_1 _09408_ (.A(_03767_),
    .B(_03768_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _09409_ (.A(net5),
    .B(net54),
    .Y(_03867_));
 sky130_fd_sc_hd__nor2_1 _09410_ (.A(_03866_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__xnor2_1 _09411_ (.A(_03765_),
    .B(_03766_),
    .Y(_03869_));
 sky130_fd_sc_hd__nand2_1 _09412_ (.A(net4),
    .B(net54),
    .Y(_03870_));
 sky130_fd_sc_hd__nor2_1 _09413_ (.A(_03869_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__xnor2_1 _09414_ (.A(_03762_),
    .B(_03764_),
    .Y(_03872_));
 sky130_fd_sc_hd__nand2_1 _09415_ (.A(net3),
    .B(net54),
    .Y(_03874_));
 sky130_fd_sc_hd__nor2_1 _09416_ (.A(_03872_),
    .B(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__xnor2_1 _09417_ (.A(_03760_),
    .B(_03761_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand2_1 _09418_ (.A(net2),
    .B(net54),
    .Y(_03877_));
 sky130_fd_sc_hd__nor2_1 _09419_ (.A(_03876_),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__xnor2_1 _09420_ (.A(_03758_),
    .B(_03759_),
    .Y(_03879_));
 sky130_fd_sc_hd__nand2_1 _09421_ (.A(net32),
    .B(net54),
    .Y(_03880_));
 sky130_fd_sc_hd__nor2_1 _09422_ (.A(_03879_),
    .B(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__xnor2_1 _09423_ (.A(_03756_),
    .B(_03757_),
    .Y(_03882_));
 sky130_fd_sc_hd__nand2_1 _09424_ (.A(net31),
    .B(net54),
    .Y(_03883_));
 sky130_fd_sc_hd__nor2_1 _09425_ (.A(_03882_),
    .B(_03883_),
    .Y(_03885_));
 sky130_fd_sc_hd__xnor2_1 _09426_ (.A(_03754_),
    .B(_03755_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand2_1 _09427_ (.A(net30),
    .B(net54),
    .Y(_03887_));
 sky130_fd_sc_hd__nor2_1 _09428_ (.A(_03886_),
    .B(_03887_),
    .Y(_03888_));
 sky130_fd_sc_hd__xnor2_1 _09429_ (.A(_03751_),
    .B(_03753_),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2_1 _09430_ (.A(net29),
    .B(net54),
    .Y(_03890_));
 sky130_fd_sc_hd__nor2_1 _09431_ (.A(_03889_),
    .B(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__xnor2_1 _09432_ (.A(_03749_),
    .B(_03750_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_1 _09433_ (.A(net28),
    .B(net54),
    .Y(_03893_));
 sky130_fd_sc_hd__nor2_1 _09434_ (.A(_03892_),
    .B(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__xnor2_1 _09435_ (.A(_03747_),
    .B(_03748_),
    .Y(_03896_));
 sky130_fd_sc_hd__nand2_1 _09436_ (.A(net27),
    .B(net54),
    .Y(_03897_));
 sky130_fd_sc_hd__nor2_1 _09437_ (.A(_03896_),
    .B(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__xnor2_1 _09438_ (.A(_03745_),
    .B(_03746_),
    .Y(_03899_));
 sky130_fd_sc_hd__nand2_1 _09439_ (.A(net26),
    .B(net54),
    .Y(_03900_));
 sky130_fd_sc_hd__nor2_1 _09440_ (.A(_03899_),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__a21o_1 _09441_ (.A1(_01470_),
    .A2(_01628_),
    .B1(_01627_),
    .X(_03902_));
 sky130_fd_sc_hd__xor2_1 _09442_ (.A(_03899_),
    .B(_03900_),
    .X(_03903_));
 sky130_fd_sc_hd__a21o_1 _09443_ (.A1(_03902_),
    .A2(_03903_),
    .B1(_03901_),
    .X(_03904_));
 sky130_fd_sc_hd__xor2_1 _09444_ (.A(_03896_),
    .B(_03897_),
    .X(_03905_));
 sky130_fd_sc_hd__a21o_1 _09445_ (.A1(_03904_),
    .A2(_03905_),
    .B1(_03898_),
    .X(_03907_));
 sky130_fd_sc_hd__xor2_1 _09446_ (.A(_03892_),
    .B(_03893_),
    .X(_03908_));
 sky130_fd_sc_hd__a21o_1 _09447_ (.A1(_03907_),
    .A2(_03908_),
    .B1(_03894_),
    .X(_03909_));
 sky130_fd_sc_hd__xor2_1 _09448_ (.A(_03889_),
    .B(_03890_),
    .X(_03910_));
 sky130_fd_sc_hd__a21o_1 _09449_ (.A1(_03909_),
    .A2(_03910_),
    .B1(_03891_),
    .X(_03911_));
 sky130_fd_sc_hd__xor2_1 _09450_ (.A(_03886_),
    .B(_03887_),
    .X(_03912_));
 sky130_fd_sc_hd__a21o_1 _09451_ (.A1(_03911_),
    .A2(_03912_),
    .B1(_03888_),
    .X(_03913_));
 sky130_fd_sc_hd__xor2_1 _09452_ (.A(_03882_),
    .B(_03883_),
    .X(_03914_));
 sky130_fd_sc_hd__a21o_1 _09453_ (.A1(_03913_),
    .A2(_03914_),
    .B1(_03885_),
    .X(_03915_));
 sky130_fd_sc_hd__xor2_1 _09454_ (.A(_03879_),
    .B(_03880_),
    .X(_03916_));
 sky130_fd_sc_hd__a21o_1 _09455_ (.A1(_03915_),
    .A2(_03916_),
    .B1(_03881_),
    .X(_03918_));
 sky130_fd_sc_hd__xor2_1 _09456_ (.A(_03876_),
    .B(_03877_),
    .X(_03919_));
 sky130_fd_sc_hd__a21o_1 _09457_ (.A1(_03918_),
    .A2(_03919_),
    .B1(_03878_),
    .X(_03920_));
 sky130_fd_sc_hd__xor2_1 _09458_ (.A(_03872_),
    .B(_03874_),
    .X(_03921_));
 sky130_fd_sc_hd__a21o_1 _09459_ (.A1(_03920_),
    .A2(_03921_),
    .B1(_03875_),
    .X(_03922_));
 sky130_fd_sc_hd__xor2_1 _09460_ (.A(_03869_),
    .B(_03870_),
    .X(_03923_));
 sky130_fd_sc_hd__a21o_1 _09461_ (.A1(_03922_),
    .A2(_03923_),
    .B1(_03871_),
    .X(_03924_));
 sky130_fd_sc_hd__xor2_1 _09462_ (.A(_03866_),
    .B(_03867_),
    .X(_03925_));
 sky130_fd_sc_hd__a21o_1 _09463_ (.A1(_03924_),
    .A2(_03925_),
    .B1(_03868_),
    .X(_03926_));
 sky130_fd_sc_hd__xor2_1 _09464_ (.A(_03863_),
    .B(_03864_),
    .X(_03927_));
 sky130_fd_sc_hd__a21o_1 _09465_ (.A1(_03926_),
    .A2(_03927_),
    .B1(_03865_),
    .X(_03929_));
 sky130_fd_sc_hd__xor2_1 _09466_ (.A(_03859_),
    .B(_03860_),
    .X(_03930_));
 sky130_fd_sc_hd__a21o_1 _09467_ (.A1(_03929_),
    .A2(_03930_),
    .B1(_03861_),
    .X(_03931_));
 sky130_fd_sc_hd__xor2_1 _09468_ (.A(_03856_),
    .B(_03857_),
    .X(_03932_));
 sky130_fd_sc_hd__a21o_1 _09469_ (.A1(_03931_),
    .A2(_03932_),
    .B1(_03858_),
    .X(_03933_));
 sky130_fd_sc_hd__xor2_1 _09470_ (.A(_03853_),
    .B(_03854_),
    .X(_03934_));
 sky130_fd_sc_hd__a21o_1 _09471_ (.A1(_03933_),
    .A2(_03934_),
    .B1(_03855_),
    .X(_03935_));
 sky130_fd_sc_hd__xor2_1 _09472_ (.A(_03849_),
    .B(_03850_),
    .X(_03936_));
 sky130_fd_sc_hd__a21o_1 _09473_ (.A1(_03935_),
    .A2(_03936_),
    .B1(_03852_),
    .X(_03937_));
 sky130_fd_sc_hd__xor2_1 _09474_ (.A(_03846_),
    .B(_03847_),
    .X(_03938_));
 sky130_fd_sc_hd__a21o_1 _09475_ (.A1(_03937_),
    .A2(_03938_),
    .B1(_03848_),
    .X(_03940_));
 sky130_fd_sc_hd__xor2_1 _09476_ (.A(_03843_),
    .B(_03844_),
    .X(_03941_));
 sky130_fd_sc_hd__a21o_1 _09477_ (.A1(_03940_),
    .A2(_03941_),
    .B1(_03845_),
    .X(_03942_));
 sky130_fd_sc_hd__xor2_1 _09478_ (.A(_03839_),
    .B(_03841_),
    .X(_03943_));
 sky130_fd_sc_hd__a21o_1 _09479_ (.A1(_03942_),
    .A2(_03943_),
    .B1(_03842_),
    .X(_03944_));
 sky130_fd_sc_hd__xor2_1 _09480_ (.A(_03836_),
    .B(_03837_),
    .X(_03945_));
 sky130_fd_sc_hd__a21o_1 _09481_ (.A1(_03944_),
    .A2(_03945_),
    .B1(_03838_),
    .X(_03946_));
 sky130_fd_sc_hd__xor2_1 _09482_ (.A(_03833_),
    .B(_03834_),
    .X(_03947_));
 sky130_fd_sc_hd__a21o_1 _09483_ (.A1(_03946_),
    .A2(_03947_),
    .B1(_03835_),
    .X(_03948_));
 sky130_fd_sc_hd__xor2_1 _09484_ (.A(_03830_),
    .B(_03831_),
    .X(_03949_));
 sky130_fd_sc_hd__a21o_1 _09485_ (.A1(_03948_),
    .A2(_03949_),
    .B1(_03832_),
    .X(_03951_));
 sky130_fd_sc_hd__xor2_1 _09486_ (.A(_03826_),
    .B(_03827_),
    .X(_03952_));
 sky130_fd_sc_hd__a21o_1 _09487_ (.A1(_03951_),
    .A2(_03952_),
    .B1(_03828_),
    .X(_03953_));
 sky130_fd_sc_hd__xor2_1 _09488_ (.A(_03823_),
    .B(_03824_),
    .X(_03954_));
 sky130_fd_sc_hd__a21o_1 _09489_ (.A1(_03953_),
    .A2(_03954_),
    .B1(_03825_),
    .X(_03955_));
 sky130_fd_sc_hd__xor2_1 _09490_ (.A(_03820_),
    .B(_03821_),
    .X(_03956_));
 sky130_fd_sc_hd__a21o_1 _09491_ (.A1(_03955_),
    .A2(_03956_),
    .B1(_03822_),
    .X(_03957_));
 sky130_fd_sc_hd__xor2_1 _09492_ (.A(_03816_),
    .B(_03817_),
    .X(_03958_));
 sky130_fd_sc_hd__a21o_1 _09493_ (.A1(_03957_),
    .A2(_03958_),
    .B1(_03819_),
    .X(_03959_));
 sky130_fd_sc_hd__xor2_1 _09494_ (.A(_03813_),
    .B(_03814_),
    .X(_03960_));
 sky130_fd_sc_hd__a21oi_1 _09495_ (.A1(_03959_),
    .A2(_03960_),
    .B1(_03815_),
    .Y(_03962_));
 sky130_fd_sc_hd__nand2_1 _09496_ (.A(net53),
    .B(net25),
    .Y(_03963_));
 sky130_fd_sc_hd__nand3_1 _09497_ (.A(_03652_),
    .B(_03803_),
    .C(_03963_),
    .Y(_03964_));
 sky130_fd_sc_hd__a21o_1 _09498_ (.A1(_03652_),
    .A2(_03803_),
    .B1(_03963_),
    .X(_03965_));
 sky130_fd_sc_hd__a211o_1 _09499_ (.A1(_03964_),
    .A2(_03965_),
    .B1(_03810_),
    .C1(_03812_),
    .X(_03966_));
 sky130_fd_sc_hd__nand2_1 _09500_ (.A(net54),
    .B(net24),
    .Y(_03967_));
 sky130_fd_sc_hd__and3_1 _09501_ (.A(net54),
    .B(net24),
    .C(_03966_),
    .X(_03968_));
 sky130_fd_sc_hd__xor2_1 _09502_ (.A(_03966_),
    .B(_03967_),
    .X(_03969_));
 sky130_fd_sc_hd__nor2_1 _09503_ (.A(_03962_),
    .B(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__xnor2_1 _09504_ (.A(_03962_),
    .B(_03969_),
    .Y(_03971_));
 sky130_fd_sc_hd__nand2_1 _09505_ (.A(net22),
    .B(net56),
    .Y(_03973_));
 sky130_fd_sc_hd__nor2_1 _09506_ (.A(_03971_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__xnor2_1 _09507_ (.A(_03959_),
    .B(_03960_),
    .Y(_03975_));
 sky130_fd_sc_hd__nand2_1 _09508_ (.A(net21),
    .B(net56),
    .Y(_03976_));
 sky130_fd_sc_hd__nor2_1 _09509_ (.A(_03975_),
    .B(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__xnor2_1 _09510_ (.A(_03957_),
    .B(_03958_),
    .Y(_03978_));
 sky130_fd_sc_hd__nand2_1 _09511_ (.A(net20),
    .B(net56),
    .Y(_03979_));
 sky130_fd_sc_hd__nor2_1 _09512_ (.A(_03978_),
    .B(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__xnor2_1 _09513_ (.A(_03955_),
    .B(_03956_),
    .Y(_03981_));
 sky130_fd_sc_hd__nand2_1 _09514_ (.A(net19),
    .B(net56),
    .Y(_03982_));
 sky130_fd_sc_hd__nor2_1 _09515_ (.A(_03981_),
    .B(_03982_),
    .Y(_03984_));
 sky130_fd_sc_hd__xnor2_1 _09516_ (.A(_03953_),
    .B(_03954_),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _09517_ (.A(net18),
    .B(net56),
    .Y(_03986_));
 sky130_fd_sc_hd__nor2_1 _09518_ (.A(_03985_),
    .B(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__xnor2_1 _09519_ (.A(_03951_),
    .B(_03952_),
    .Y(_03988_));
 sky130_fd_sc_hd__nand2_1 _09520_ (.A(net17),
    .B(net56),
    .Y(_03989_));
 sky130_fd_sc_hd__nor2_1 _09521_ (.A(_03988_),
    .B(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__xnor2_1 _09522_ (.A(_03948_),
    .B(_03949_),
    .Y(_03991_));
 sky130_fd_sc_hd__nand2_1 _09523_ (.A(net16),
    .B(net56),
    .Y(_03992_));
 sky130_fd_sc_hd__nor2_1 _09524_ (.A(_03991_),
    .B(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__xnor2_1 _09525_ (.A(_03946_),
    .B(_03947_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand2_1 _09526_ (.A(net15),
    .B(net56),
    .Y(_03996_));
 sky130_fd_sc_hd__nor2_1 _09527_ (.A(_03995_),
    .B(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__xnor2_1 _09528_ (.A(_03944_),
    .B(_03945_),
    .Y(_03998_));
 sky130_fd_sc_hd__nand2_1 _09529_ (.A(net14),
    .B(net56),
    .Y(_03999_));
 sky130_fd_sc_hd__nor2_1 _09530_ (.A(_03998_),
    .B(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__xnor2_1 _09531_ (.A(_03942_),
    .B(_03943_),
    .Y(_04001_));
 sky130_fd_sc_hd__nand2_1 _09532_ (.A(net13),
    .B(net56),
    .Y(_04002_));
 sky130_fd_sc_hd__nor2_1 _09533_ (.A(_04001_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__xnor2_1 _09534_ (.A(_03940_),
    .B(_03941_),
    .Y(_04004_));
 sky130_fd_sc_hd__nand2_1 _09535_ (.A(net11),
    .B(net56),
    .Y(_04006_));
 sky130_fd_sc_hd__nor2_1 _09536_ (.A(_04004_),
    .B(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__xnor2_1 _09537_ (.A(_03937_),
    .B(_03938_),
    .Y(_04008_));
 sky130_fd_sc_hd__nand2_1 _09538_ (.A(net10),
    .B(net56),
    .Y(_04009_));
 sky130_fd_sc_hd__nor2_1 _09539_ (.A(_04008_),
    .B(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__xnor2_1 _09540_ (.A(_03935_),
    .B(_03936_),
    .Y(_04011_));
 sky130_fd_sc_hd__nand2_1 _09541_ (.A(net9),
    .B(net56),
    .Y(_04012_));
 sky130_fd_sc_hd__nor2_1 _09542_ (.A(_04011_),
    .B(_04012_),
    .Y(_04013_));
 sky130_fd_sc_hd__xnor2_1 _09543_ (.A(_03933_),
    .B(_03934_),
    .Y(_04014_));
 sky130_fd_sc_hd__nand2_1 _09544_ (.A(net8),
    .B(net56),
    .Y(_04015_));
 sky130_fd_sc_hd__nor2_1 _09545_ (.A(_04014_),
    .B(_04015_),
    .Y(_04017_));
 sky130_fd_sc_hd__xnor2_1 _09546_ (.A(_03931_),
    .B(_03932_),
    .Y(_04018_));
 sky130_fd_sc_hd__nand2_1 _09547_ (.A(net7),
    .B(net56),
    .Y(_04019_));
 sky130_fd_sc_hd__nor2_1 _09548_ (.A(_04018_),
    .B(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__xnor2_1 _09549_ (.A(_03929_),
    .B(_03930_),
    .Y(_04021_));
 sky130_fd_sc_hd__nand2_1 _09550_ (.A(net6),
    .B(net56),
    .Y(_04022_));
 sky130_fd_sc_hd__nor2_1 _09551_ (.A(_04021_),
    .B(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__xnor2_1 _09552_ (.A(_03926_),
    .B(_03927_),
    .Y(_04024_));
 sky130_fd_sc_hd__nand2_1 _09553_ (.A(net5),
    .B(net56),
    .Y(_04025_));
 sky130_fd_sc_hd__nor2_1 _09554_ (.A(_04024_),
    .B(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__xnor2_1 _09555_ (.A(_03924_),
    .B(_03925_),
    .Y(_04028_));
 sky130_fd_sc_hd__nand2_1 _09556_ (.A(net4),
    .B(net56),
    .Y(_04029_));
 sky130_fd_sc_hd__nor2_1 _09557_ (.A(_04028_),
    .B(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__xnor2_1 _09558_ (.A(_03922_),
    .B(_03923_),
    .Y(_04031_));
 sky130_fd_sc_hd__nand2_1 _09559_ (.A(net3),
    .B(net56),
    .Y(_04032_));
 sky130_fd_sc_hd__nor2_1 _09560_ (.A(_04031_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__xnor2_1 _09561_ (.A(_03920_),
    .B(_03921_),
    .Y(_04034_));
 sky130_fd_sc_hd__nand2_1 _09562_ (.A(net2),
    .B(net56),
    .Y(_04035_));
 sky130_fd_sc_hd__nor2_1 _09563_ (.A(_04034_),
    .B(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__xnor2_1 _09564_ (.A(_03918_),
    .B(_03919_),
    .Y(_04037_));
 sky130_fd_sc_hd__nand2_1 _09565_ (.A(net32),
    .B(net56),
    .Y(_04039_));
 sky130_fd_sc_hd__nor2_1 _09566_ (.A(_04037_),
    .B(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__xnor2_1 _09567_ (.A(_03915_),
    .B(_03916_),
    .Y(_04041_));
 sky130_fd_sc_hd__nand2_1 _09568_ (.A(net31),
    .B(net56),
    .Y(_04042_));
 sky130_fd_sc_hd__nor2_1 _09569_ (.A(_04041_),
    .B(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__xnor2_1 _09570_ (.A(_03913_),
    .B(_03914_),
    .Y(_04044_));
 sky130_fd_sc_hd__nand2_1 _09571_ (.A(net30),
    .B(net56),
    .Y(_04045_));
 sky130_fd_sc_hd__nor2_1 _09572_ (.A(_04044_),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__xnor2_1 _09573_ (.A(_03911_),
    .B(_03912_),
    .Y(_04047_));
 sky130_fd_sc_hd__nand2_1 _09574_ (.A(net29),
    .B(net56),
    .Y(_04048_));
 sky130_fd_sc_hd__nor2_1 _09575_ (.A(_04047_),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__xnor2_1 _09576_ (.A(_03909_),
    .B(_03910_),
    .Y(_04050_));
 sky130_fd_sc_hd__nand2_1 _09577_ (.A(net28),
    .B(net56),
    .Y(_04051_));
 sky130_fd_sc_hd__nor2_1 _09578_ (.A(_04050_),
    .B(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__xnor2_1 _09579_ (.A(_03907_),
    .B(_03908_),
    .Y(_04053_));
 sky130_fd_sc_hd__nand2_1 _09580_ (.A(net27),
    .B(net56),
    .Y(_04054_));
 sky130_fd_sc_hd__nor2_1 _09581_ (.A(_04053_),
    .B(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__xnor2_1 _09582_ (.A(_03904_),
    .B(_03905_),
    .Y(_04056_));
 sky130_fd_sc_hd__nand2_1 _09583_ (.A(net26),
    .B(net56),
    .Y(_04057_));
 sky130_fd_sc_hd__nor2_1 _09584_ (.A(_04056_),
    .B(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__xnor2_1 _09585_ (.A(_03902_),
    .B(_03903_),
    .Y(_04060_));
 sky130_fd_sc_hd__nand2_1 _09586_ (.A(net23),
    .B(net56),
    .Y(_04061_));
 sky130_fd_sc_hd__nor2_1 _09587_ (.A(_04060_),
    .B(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__a21o_1 _09588_ (.A1(_01467_),
    .A2(_01632_),
    .B1(_01631_),
    .X(_04063_));
 sky130_fd_sc_hd__xor2_1 _09589_ (.A(_04060_),
    .B(_04061_),
    .X(_04064_));
 sky130_fd_sc_hd__a21o_1 _09590_ (.A1(_04063_),
    .A2(_04064_),
    .B1(_04062_),
    .X(_04065_));
 sky130_fd_sc_hd__xor2_1 _09591_ (.A(_04056_),
    .B(_04057_),
    .X(_04066_));
 sky130_fd_sc_hd__a21o_1 _09592_ (.A1(_04065_),
    .A2(_04066_),
    .B1(_04058_),
    .X(_04067_));
 sky130_fd_sc_hd__xor2_1 _09593_ (.A(_04053_),
    .B(_04054_),
    .X(_04068_));
 sky130_fd_sc_hd__a21o_1 _09594_ (.A1(_04067_),
    .A2(_04068_),
    .B1(_04055_),
    .X(_04069_));
 sky130_fd_sc_hd__xor2_1 _09595_ (.A(_04050_),
    .B(_04051_),
    .X(_04071_));
 sky130_fd_sc_hd__a21o_1 _09596_ (.A1(_04069_),
    .A2(_04071_),
    .B1(_04052_),
    .X(_04072_));
 sky130_fd_sc_hd__xor2_1 _09597_ (.A(_04047_),
    .B(_04048_),
    .X(_04073_));
 sky130_fd_sc_hd__a21o_1 _09598_ (.A1(_04072_),
    .A2(_04073_),
    .B1(_04049_),
    .X(_04074_));
 sky130_fd_sc_hd__xor2_1 _09599_ (.A(_04044_),
    .B(_04045_),
    .X(_04075_));
 sky130_fd_sc_hd__a21o_1 _09600_ (.A1(_04074_),
    .A2(_04075_),
    .B1(_04046_),
    .X(_04076_));
 sky130_fd_sc_hd__xor2_1 _09601_ (.A(_04041_),
    .B(_04042_),
    .X(_04077_));
 sky130_fd_sc_hd__a21o_1 _09602_ (.A1(_04076_),
    .A2(_04077_),
    .B1(_04043_),
    .X(_04078_));
 sky130_fd_sc_hd__xor2_1 _09603_ (.A(_04037_),
    .B(_04039_),
    .X(_04079_));
 sky130_fd_sc_hd__a21o_1 _09604_ (.A1(_04078_),
    .A2(_04079_),
    .B1(_04040_),
    .X(_04080_));
 sky130_fd_sc_hd__xor2_1 _09605_ (.A(_04034_),
    .B(_04035_),
    .X(_04082_));
 sky130_fd_sc_hd__a21o_1 _09606_ (.A1(_04080_),
    .A2(_04082_),
    .B1(_04036_),
    .X(_04083_));
 sky130_fd_sc_hd__xor2_1 _09607_ (.A(_04031_),
    .B(_04032_),
    .X(_04084_));
 sky130_fd_sc_hd__a21o_1 _09608_ (.A1(_04083_),
    .A2(_04084_),
    .B1(_04033_),
    .X(_04085_));
 sky130_fd_sc_hd__xor2_1 _09609_ (.A(_04028_),
    .B(_04029_),
    .X(_04086_));
 sky130_fd_sc_hd__a21o_1 _09610_ (.A1(_04085_),
    .A2(_04086_),
    .B1(_04030_),
    .X(_04087_));
 sky130_fd_sc_hd__xor2_1 _09611_ (.A(_04024_),
    .B(_04025_),
    .X(_04088_));
 sky130_fd_sc_hd__a21o_1 _09612_ (.A1(_04087_),
    .A2(_04088_),
    .B1(_04026_),
    .X(_04089_));
 sky130_fd_sc_hd__xor2_1 _09613_ (.A(_04021_),
    .B(_04022_),
    .X(_04090_));
 sky130_fd_sc_hd__a21o_1 _09614_ (.A1(_04089_),
    .A2(_04090_),
    .B1(_04023_),
    .X(_04091_));
 sky130_fd_sc_hd__xor2_1 _09615_ (.A(_04018_),
    .B(_04019_),
    .X(_04093_));
 sky130_fd_sc_hd__a21o_1 _09616_ (.A1(_04091_),
    .A2(_04093_),
    .B1(_04020_),
    .X(_04094_));
 sky130_fd_sc_hd__xor2_1 _09617_ (.A(_04014_),
    .B(_04015_),
    .X(_04095_));
 sky130_fd_sc_hd__a21o_1 _09618_ (.A1(_04094_),
    .A2(_04095_),
    .B1(_04017_),
    .X(_04096_));
 sky130_fd_sc_hd__xor2_1 _09619_ (.A(_04011_),
    .B(_04012_),
    .X(_04097_));
 sky130_fd_sc_hd__a21o_1 _09620_ (.A1(_04096_),
    .A2(_04097_),
    .B1(_04013_),
    .X(_04098_));
 sky130_fd_sc_hd__xor2_1 _09621_ (.A(_04008_),
    .B(_04009_),
    .X(_04099_));
 sky130_fd_sc_hd__a21o_1 _09622_ (.A1(_04098_),
    .A2(_04099_),
    .B1(_04010_),
    .X(_04100_));
 sky130_fd_sc_hd__xor2_1 _09623_ (.A(_04004_),
    .B(_04006_),
    .X(_04101_));
 sky130_fd_sc_hd__a21o_1 _09624_ (.A1(_04100_),
    .A2(_04101_),
    .B1(_04007_),
    .X(_04102_));
 sky130_fd_sc_hd__xor2_1 _09625_ (.A(_04001_),
    .B(_04002_),
    .X(_04104_));
 sky130_fd_sc_hd__a21o_1 _09626_ (.A1(_04102_),
    .A2(_04104_),
    .B1(_04003_),
    .X(_04105_));
 sky130_fd_sc_hd__xor2_1 _09627_ (.A(_03998_),
    .B(_03999_),
    .X(_04106_));
 sky130_fd_sc_hd__a21o_1 _09628_ (.A1(_04105_),
    .A2(_04106_),
    .B1(_04000_),
    .X(_04107_));
 sky130_fd_sc_hd__xor2_1 _09629_ (.A(_03995_),
    .B(_03996_),
    .X(_04108_));
 sky130_fd_sc_hd__a21o_1 _09630_ (.A1(_04107_),
    .A2(_04108_),
    .B1(_03997_),
    .X(_04109_));
 sky130_fd_sc_hd__xor2_1 _09631_ (.A(_03991_),
    .B(_03992_),
    .X(_04110_));
 sky130_fd_sc_hd__a21o_1 _09632_ (.A1(_04109_),
    .A2(_04110_),
    .B1(_03993_),
    .X(_04111_));
 sky130_fd_sc_hd__xor2_1 _09633_ (.A(_03988_),
    .B(_03989_),
    .X(_04112_));
 sky130_fd_sc_hd__a21o_1 _09634_ (.A1(_04111_),
    .A2(_04112_),
    .B1(_03990_),
    .X(_04113_));
 sky130_fd_sc_hd__xor2_1 _09635_ (.A(_03985_),
    .B(_03986_),
    .X(_04115_));
 sky130_fd_sc_hd__a21o_1 _09636_ (.A1(_04113_),
    .A2(_04115_),
    .B1(_03987_),
    .X(_04116_));
 sky130_fd_sc_hd__xor2_1 _09637_ (.A(_03981_),
    .B(_03982_),
    .X(_04117_));
 sky130_fd_sc_hd__a21o_1 _09638_ (.A1(_04116_),
    .A2(_04117_),
    .B1(_03984_),
    .X(_04118_));
 sky130_fd_sc_hd__xor2_1 _09639_ (.A(_03978_),
    .B(_03979_),
    .X(_04119_));
 sky130_fd_sc_hd__a21o_1 _09640_ (.A1(_04118_),
    .A2(_04119_),
    .B1(_03980_),
    .X(_04120_));
 sky130_fd_sc_hd__xor2_1 _09641_ (.A(_03975_),
    .B(_03976_),
    .X(_04121_));
 sky130_fd_sc_hd__a21o_1 _09642_ (.A1(_04120_),
    .A2(_04121_),
    .B1(_03977_),
    .X(_04122_));
 sky130_fd_sc_hd__xor2_1 _09643_ (.A(_03971_),
    .B(_03973_),
    .X(_04123_));
 sky130_fd_sc_hd__a21oi_1 _09644_ (.A1(_04122_),
    .A2(_04123_),
    .B1(_03974_),
    .Y(_04124_));
 sky130_fd_sc_hd__nand2_1 _09645_ (.A(net54),
    .B(net25),
    .Y(_04126_));
 sky130_fd_sc_hd__nand2b_1 _09646_ (.A_N(_03964_),
    .B(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__and3_1 _09647_ (.A(net54),
    .B(net25),
    .C(_03964_),
    .X(_04128_));
 sky130_fd_sc_hd__inv_2 _09648_ (.A(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__a211o_1 _09649_ (.A1(_04127_),
    .A2(_04129_),
    .B1(_03968_),
    .C1(_03970_),
    .X(_04130_));
 sky130_fd_sc_hd__and2_1 _09650_ (.A(net24),
    .B(net56),
    .X(_04131_));
 sky130_fd_sc_hd__nand2_1 _09651_ (.A(_04130_),
    .B(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__xnor2_1 _09652_ (.A(_04130_),
    .B(_04131_),
    .Y(_04133_));
 sky130_fd_sc_hd__xnor2_1 _09653_ (.A(_04124_),
    .B(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__or2_1 _09654_ (.A(net12),
    .B(net1),
    .X(_04135_));
 sky130_fd_sc_hd__or2_1 _09655_ (.A(net23),
    .B(_04135_),
    .X(_04137_));
 sky130_fd_sc_hd__or2_1 _09656_ (.A(net26),
    .B(_04137_),
    .X(_04138_));
 sky130_fd_sc_hd__or2_1 _09657_ (.A(net27),
    .B(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__or2_1 _09658_ (.A(net28),
    .B(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__or2_1 _09659_ (.A(net29),
    .B(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__or2_1 _09660_ (.A(net30),
    .B(_04141_),
    .X(_04142_));
 sky130_fd_sc_hd__or2_1 _09661_ (.A(net31),
    .B(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__or2_1 _09662_ (.A(net32),
    .B(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__or2_1 _09663_ (.A(net2),
    .B(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__or2_1 _09664_ (.A(net3),
    .B(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__or2_1 _09665_ (.A(net4),
    .B(_04146_),
    .X(_04148_));
 sky130_fd_sc_hd__or2_1 _09666_ (.A(net5),
    .B(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__or2_1 _09667_ (.A(net6),
    .B(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__or2_1 _09668_ (.A(net7),
    .B(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__or2_1 _09669_ (.A(net8),
    .B(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__or2_1 _09670_ (.A(net9),
    .B(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__or2_1 _09671_ (.A(net10),
    .B(_04153_),
    .X(_04154_));
 sky130_fd_sc_hd__or2_1 _09672_ (.A(net11),
    .B(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__or2_1 _09673_ (.A(net13),
    .B(_04155_),
    .X(_04156_));
 sky130_fd_sc_hd__or2_1 _09674_ (.A(net14),
    .B(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__or2_1 _09675_ (.A(net15),
    .B(_04157_),
    .X(_04159_));
 sky130_fd_sc_hd__or2_1 _09676_ (.A(net16),
    .B(_04159_),
    .X(_04160_));
 sky130_fd_sc_hd__or2_1 _09677_ (.A(net17),
    .B(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__or2_1 _09678_ (.A(net18),
    .B(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__or2_1 _09679_ (.A(net19),
    .B(_04162_),
    .X(_04163_));
 sky130_fd_sc_hd__or2_1 _09680_ (.A(net20),
    .B(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__or2_1 _09681_ (.A(net21),
    .B(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__nand2_1 _09682_ (.A(net22),
    .B(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__or2_1 _09683_ (.A(net22),
    .B(_04165_),
    .X(_04167_));
 sky130_fd_sc_hd__and3_1 _09684_ (.A(net57),
    .B(_04166_),
    .C(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__inv_2 _09685_ (.A(_04168_),
    .Y(_04170_));
 sky130_fd_sc_hd__nor2_1 _09686_ (.A(_04134_),
    .B(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__xnor2_1 _09687_ (.A(_04122_),
    .B(_04123_),
    .Y(_04172_));
 sky130_fd_sc_hd__nand2_1 _09688_ (.A(net21),
    .B(_04164_),
    .Y(_04173_));
 sky130_fd_sc_hd__and3_1 _09689_ (.A(net57),
    .B(_04165_),
    .C(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__inv_2 _09690_ (.A(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__nor2_1 _09691_ (.A(_04172_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__xnor2_1 _09692_ (.A(_04120_),
    .B(_04121_),
    .Y(_04177_));
 sky130_fd_sc_hd__nand2_1 _09693_ (.A(net20),
    .B(_04163_),
    .Y(_04178_));
 sky130_fd_sc_hd__and3_1 _09694_ (.A(net57),
    .B(_04164_),
    .C(_04178_),
    .X(_04179_));
 sky130_fd_sc_hd__inv_2 _09695_ (.A(_04179_),
    .Y(_04181_));
 sky130_fd_sc_hd__nor2_1 _09696_ (.A(_04177_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__xnor2_1 _09697_ (.A(_04118_),
    .B(_04119_),
    .Y(_04183_));
 sky130_fd_sc_hd__nand2_1 _09698_ (.A(net19),
    .B(_04162_),
    .Y(_04184_));
 sky130_fd_sc_hd__and3_1 _09699_ (.A(net57),
    .B(_04163_),
    .C(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__inv_2 _09700_ (.A(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__nor2_1 _09701_ (.A(_04183_),
    .B(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__xnor2_1 _09702_ (.A(_04116_),
    .B(_04117_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand2_1 _09703_ (.A(net18),
    .B(_04161_),
    .Y(_04189_));
 sky130_fd_sc_hd__and3_1 _09704_ (.A(net57),
    .B(_04162_),
    .C(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__inv_2 _09705_ (.A(_04190_),
    .Y(_04192_));
 sky130_fd_sc_hd__nor2_1 _09706_ (.A(_04188_),
    .B(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__xnor2_1 _09707_ (.A(_04113_),
    .B(_04115_),
    .Y(_04194_));
 sky130_fd_sc_hd__nand2_1 _09708_ (.A(net17),
    .B(_04160_),
    .Y(_04195_));
 sky130_fd_sc_hd__and3_1 _09709_ (.A(net57),
    .B(_04161_),
    .C(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__inv_2 _09710_ (.A(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__nor2_1 _09711_ (.A(_04194_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__xnor2_1 _09712_ (.A(_04111_),
    .B(_04112_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand2_1 _09713_ (.A(net16),
    .B(_04159_),
    .Y(_04200_));
 sky130_fd_sc_hd__and3_1 _09714_ (.A(net57),
    .B(_04160_),
    .C(_04200_),
    .X(_04201_));
 sky130_fd_sc_hd__inv_2 _09715_ (.A(_04201_),
    .Y(_04203_));
 sky130_fd_sc_hd__nor2_1 _09716_ (.A(_04199_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__xnor2_1 _09717_ (.A(_04109_),
    .B(_04110_),
    .Y(_04205_));
 sky130_fd_sc_hd__nand2_1 _09718_ (.A(net15),
    .B(_04157_),
    .Y(_04206_));
 sky130_fd_sc_hd__and3_1 _09719_ (.A(net57),
    .B(_04159_),
    .C(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__inv_2 _09720_ (.A(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__nor2_1 _09721_ (.A(_04205_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__xnor2_1 _09722_ (.A(_04107_),
    .B(_04108_),
    .Y(_04210_));
 sky130_fd_sc_hd__nand2_1 _09723_ (.A(net14),
    .B(_04156_),
    .Y(_04211_));
 sky130_fd_sc_hd__and3_1 _09724_ (.A(net57),
    .B(_04157_),
    .C(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__inv_2 _09725_ (.A(_04212_),
    .Y(_04214_));
 sky130_fd_sc_hd__nor2_1 _09726_ (.A(_04210_),
    .B(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__xnor2_1 _09727_ (.A(_04105_),
    .B(_04106_),
    .Y(_04216_));
 sky130_fd_sc_hd__nand2_1 _09728_ (.A(net13),
    .B(_04155_),
    .Y(_04217_));
 sky130_fd_sc_hd__and3_1 _09729_ (.A(net57),
    .B(_04156_),
    .C(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__inv_2 _09730_ (.A(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__nor2_1 _09731_ (.A(_04216_),
    .B(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__xnor2_1 _09732_ (.A(_04102_),
    .B(_04104_),
    .Y(_04221_));
 sky130_fd_sc_hd__nand2_1 _09733_ (.A(net11),
    .B(_04154_),
    .Y(_04222_));
 sky130_fd_sc_hd__and3_1 _09734_ (.A(net57),
    .B(_04155_),
    .C(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__inv_2 _09735_ (.A(_04223_),
    .Y(_04225_));
 sky130_fd_sc_hd__nor2_1 _09736_ (.A(_04221_),
    .B(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__xnor2_1 _09737_ (.A(_04100_),
    .B(_04101_),
    .Y(_04227_));
 sky130_fd_sc_hd__nand2_1 _09738_ (.A(net10),
    .B(_04153_),
    .Y(_04228_));
 sky130_fd_sc_hd__and3_1 _09739_ (.A(net57),
    .B(_04154_),
    .C(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__inv_2 _09740_ (.A(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__nor2_1 _09741_ (.A(_04227_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__xnor2_1 _09742_ (.A(_04098_),
    .B(_04099_),
    .Y(_04232_));
 sky130_fd_sc_hd__nand2_1 _09743_ (.A(net9),
    .B(_04152_),
    .Y(_04233_));
 sky130_fd_sc_hd__and3_1 _09744_ (.A(net57),
    .B(_04153_),
    .C(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__inv_2 _09745_ (.A(_04234_),
    .Y(_04236_));
 sky130_fd_sc_hd__nor2_1 _09746_ (.A(_04232_),
    .B(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__xnor2_1 _09747_ (.A(_04096_),
    .B(_04097_),
    .Y(_04238_));
 sky130_fd_sc_hd__nand2_1 _09748_ (.A(net8),
    .B(_04151_),
    .Y(_04239_));
 sky130_fd_sc_hd__and3_1 _09749_ (.A(net57),
    .B(_04152_),
    .C(_04239_),
    .X(_04240_));
 sky130_fd_sc_hd__inv_2 _09750_ (.A(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__nor2_1 _09751_ (.A(_04238_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__xnor2_1 _09752_ (.A(_04094_),
    .B(_04095_),
    .Y(_04243_));
 sky130_fd_sc_hd__nand2_1 _09753_ (.A(net7),
    .B(_04150_),
    .Y(_04244_));
 sky130_fd_sc_hd__and3_1 _09754_ (.A(net57),
    .B(_04151_),
    .C(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__inv_2 _09755_ (.A(_04245_),
    .Y(_04247_));
 sky130_fd_sc_hd__nor2_1 _09756_ (.A(_04243_),
    .B(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__xnor2_1 _09757_ (.A(_04091_),
    .B(_04093_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand2_1 _09758_ (.A(net6),
    .B(_04149_),
    .Y(_04250_));
 sky130_fd_sc_hd__and3_1 _09759_ (.A(net57),
    .B(_04150_),
    .C(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__inv_2 _09760_ (.A(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__nor2_1 _09761_ (.A(_04249_),
    .B(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__xnor2_1 _09762_ (.A(_04089_),
    .B(_04090_),
    .Y(_04254_));
 sky130_fd_sc_hd__nand2_1 _09763_ (.A(net5),
    .B(_04148_),
    .Y(_04255_));
 sky130_fd_sc_hd__and3_1 _09764_ (.A(net57),
    .B(_04149_),
    .C(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__inv_2 _09765_ (.A(_04256_),
    .Y(_04258_));
 sky130_fd_sc_hd__nor2_1 _09766_ (.A(_04254_),
    .B(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__xnor2_1 _09767_ (.A(_04087_),
    .B(_04088_),
    .Y(_04260_));
 sky130_fd_sc_hd__nand2_1 _09768_ (.A(net4),
    .B(_04146_),
    .Y(_04261_));
 sky130_fd_sc_hd__and3_1 _09769_ (.A(net57),
    .B(_04148_),
    .C(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__inv_2 _09770_ (.A(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__nor2_1 _09771_ (.A(_04260_),
    .B(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__xnor2_1 _09772_ (.A(_04085_),
    .B(_04086_),
    .Y(_04265_));
 sky130_fd_sc_hd__nand2_1 _09773_ (.A(net3),
    .B(_04145_),
    .Y(_04266_));
 sky130_fd_sc_hd__and3_1 _09774_ (.A(net57),
    .B(_04146_),
    .C(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__inv_2 _09775_ (.A(_04267_),
    .Y(_04269_));
 sky130_fd_sc_hd__nor2_1 _09776_ (.A(_04265_),
    .B(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__xnor2_1 _09777_ (.A(_04083_),
    .B(_04084_),
    .Y(_04271_));
 sky130_fd_sc_hd__nand2_1 _09778_ (.A(net2),
    .B(_04144_),
    .Y(_04272_));
 sky130_fd_sc_hd__and3_1 _09779_ (.A(net57),
    .B(_04145_),
    .C(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__inv_2 _09780_ (.A(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__nor2_1 _09781_ (.A(_04271_),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__xnor2_1 _09782_ (.A(_04080_),
    .B(_04082_),
    .Y(_04276_));
 sky130_fd_sc_hd__nand2_1 _09783_ (.A(net32),
    .B(_04143_),
    .Y(_04277_));
 sky130_fd_sc_hd__and3_1 _09784_ (.A(net57),
    .B(_04144_),
    .C(_04277_),
    .X(_04278_));
 sky130_fd_sc_hd__inv_2 _09785_ (.A(_04278_),
    .Y(_04280_));
 sky130_fd_sc_hd__nor2_1 _09786_ (.A(_04276_),
    .B(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__xnor2_1 _09787_ (.A(_04078_),
    .B(_04079_),
    .Y(_04282_));
 sky130_fd_sc_hd__nand2_1 _09788_ (.A(net31),
    .B(_04142_),
    .Y(_04283_));
 sky130_fd_sc_hd__and3_1 _09789_ (.A(net57),
    .B(_04143_),
    .C(_04283_),
    .X(_04284_));
 sky130_fd_sc_hd__inv_2 _09790_ (.A(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__nor2_1 _09791_ (.A(_04282_),
    .B(_04285_),
    .Y(_04286_));
 sky130_fd_sc_hd__xnor2_1 _09792_ (.A(_04076_),
    .B(_04077_),
    .Y(_04287_));
 sky130_fd_sc_hd__nand2_1 _09793_ (.A(net30),
    .B(_04141_),
    .Y(_04288_));
 sky130_fd_sc_hd__and3_1 _09794_ (.A(net57),
    .B(_04142_),
    .C(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__inv_2 _09795_ (.A(_04289_),
    .Y(_04291_));
 sky130_fd_sc_hd__nor2_1 _09796_ (.A(_04287_),
    .B(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__xnor2_1 _09797_ (.A(_04074_),
    .B(_04075_),
    .Y(_04293_));
 sky130_fd_sc_hd__nand2_1 _09798_ (.A(net29),
    .B(_04140_),
    .Y(_04294_));
 sky130_fd_sc_hd__and3_1 _09799_ (.A(net57),
    .B(_04141_),
    .C(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__inv_2 _09800_ (.A(_04295_),
    .Y(_04296_));
 sky130_fd_sc_hd__nor2_1 _09801_ (.A(_04293_),
    .B(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__xnor2_1 _09802_ (.A(_04072_),
    .B(_04073_),
    .Y(_04298_));
 sky130_fd_sc_hd__nand2_1 _09803_ (.A(net28),
    .B(_04139_),
    .Y(_04299_));
 sky130_fd_sc_hd__and3_1 _09804_ (.A(net57),
    .B(_04140_),
    .C(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__inv_2 _09805_ (.A(_04300_),
    .Y(_04302_));
 sky130_fd_sc_hd__nor2_1 _09806_ (.A(_04298_),
    .B(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__xnor2_1 _09807_ (.A(_04069_),
    .B(_04071_),
    .Y(_04304_));
 sky130_fd_sc_hd__nand2_1 _09808_ (.A(net27),
    .B(_04138_),
    .Y(_04305_));
 sky130_fd_sc_hd__and3_1 _09809_ (.A(net57),
    .B(_04139_),
    .C(_04305_),
    .X(_04306_));
 sky130_fd_sc_hd__inv_2 _09810_ (.A(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__nor2_1 _09811_ (.A(_04304_),
    .B(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__xnor2_1 _09812_ (.A(_04067_),
    .B(_04068_),
    .Y(_04309_));
 sky130_fd_sc_hd__nand2_1 _09813_ (.A(net26),
    .B(_04137_),
    .Y(_04310_));
 sky130_fd_sc_hd__and3_1 _09814_ (.A(net57),
    .B(_04138_),
    .C(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__inv_2 _09815_ (.A(_04311_),
    .Y(_04313_));
 sky130_fd_sc_hd__nor2_1 _09816_ (.A(_04309_),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__xor2_1 _09817_ (.A(_04065_),
    .B(_04066_),
    .X(_04315_));
 sky130_fd_sc_hd__nand2_1 _09818_ (.A(net23),
    .B(_04135_),
    .Y(_04316_));
 sky130_fd_sc_hd__and3_1 _09819_ (.A(net57),
    .B(_04137_),
    .C(_04316_),
    .X(_04317_));
 sky130_fd_sc_hd__and2_1 _09820_ (.A(_04315_),
    .B(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__xnor2_1 _09821_ (.A(_04063_),
    .B(_04064_),
    .Y(_04319_));
 sky130_fd_sc_hd__and3_1 _09822_ (.A(net57),
    .B(_00395_),
    .C(_04135_),
    .X(_04320_));
 sky130_fd_sc_hd__and2b_1 _09823_ (.A_N(_04319_),
    .B(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__xnor2_1 _09824_ (.A(_04319_),
    .B(_04320_),
    .Y(_04322_));
 sky130_fd_sc_hd__a21o_1 _09825_ (.A1(_01634_),
    .A2(_04322_),
    .B1(_04321_),
    .X(_04324_));
 sky130_fd_sc_hd__xor2_1 _09826_ (.A(_04315_),
    .B(_04317_),
    .X(_04325_));
 sky130_fd_sc_hd__a21o_1 _09827_ (.A1(_04324_),
    .A2(_04325_),
    .B1(_04318_),
    .X(_04326_));
 sky130_fd_sc_hd__nand2_1 _09828_ (.A(_04309_),
    .B(_04313_),
    .Y(_04327_));
 sky130_fd_sc_hd__nand2b_1 _09829_ (.A_N(_04314_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__a21o_1 _09830_ (.A1(_04326_),
    .A2(_04327_),
    .B1(_04314_),
    .X(_04329_));
 sky130_fd_sc_hd__nand2_1 _09831_ (.A(_04304_),
    .B(_04307_),
    .Y(_04330_));
 sky130_fd_sc_hd__nand2b_1 _09832_ (.A_N(_04308_),
    .B(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__a21o_1 _09833_ (.A1(_04329_),
    .A2(_04330_),
    .B1(_04308_),
    .X(_04332_));
 sky130_fd_sc_hd__nand2_1 _09834_ (.A(_04298_),
    .B(_04302_),
    .Y(_04333_));
 sky130_fd_sc_hd__nand2b_1 _09835_ (.A_N(_04303_),
    .B(_04333_),
    .Y(_04335_));
 sky130_fd_sc_hd__a21o_1 _09836_ (.A1(_04332_),
    .A2(_04333_),
    .B1(_04303_),
    .X(_04336_));
 sky130_fd_sc_hd__nand2_1 _09837_ (.A(_04293_),
    .B(_04296_),
    .Y(_04337_));
 sky130_fd_sc_hd__nand2b_1 _09838_ (.A_N(_04297_),
    .B(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__a21o_1 _09839_ (.A1(_04336_),
    .A2(_04337_),
    .B1(_04297_),
    .X(_04339_));
 sky130_fd_sc_hd__nand2_1 _09840_ (.A(_04287_),
    .B(_04291_),
    .Y(_04340_));
 sky130_fd_sc_hd__nand2b_1 _09841_ (.A_N(_04292_),
    .B(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__a21o_1 _09842_ (.A1(_04339_),
    .A2(_04340_),
    .B1(_04292_),
    .X(_04342_));
 sky130_fd_sc_hd__nand2_1 _09843_ (.A(_04282_),
    .B(_04285_),
    .Y(_04343_));
 sky130_fd_sc_hd__nand2b_1 _09844_ (.A_N(_04286_),
    .B(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__a21o_1 _09845_ (.A1(_04342_),
    .A2(_04343_),
    .B1(_04286_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _09846_ (.A(_04276_),
    .B(_04280_),
    .Y(_04347_));
 sky130_fd_sc_hd__nand2b_1 _09847_ (.A_N(_04281_),
    .B(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__a21o_1 _09848_ (.A1(_04346_),
    .A2(_04347_),
    .B1(_04281_),
    .X(_04349_));
 sky130_fd_sc_hd__nand2_1 _09849_ (.A(_04271_),
    .B(_04274_),
    .Y(_04350_));
 sky130_fd_sc_hd__nand2b_1 _09850_ (.A_N(_04275_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__a21o_1 _09851_ (.A1(_04349_),
    .A2(_04350_),
    .B1(_04275_),
    .X(_04352_));
 sky130_fd_sc_hd__nand2_1 _09852_ (.A(_04265_),
    .B(_04269_),
    .Y(_04353_));
 sky130_fd_sc_hd__nand2b_1 _09853_ (.A_N(_04270_),
    .B(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__a21o_1 _09854_ (.A1(_04352_),
    .A2(_04353_),
    .B1(_04270_),
    .X(_04355_));
 sky130_fd_sc_hd__nand2_1 _09855_ (.A(_04260_),
    .B(_04263_),
    .Y(_04357_));
 sky130_fd_sc_hd__nand2b_1 _09856_ (.A_N(_04264_),
    .B(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__a21o_1 _09857_ (.A1(_04355_),
    .A2(_04357_),
    .B1(_04264_),
    .X(_04359_));
 sky130_fd_sc_hd__nand2_1 _09858_ (.A(_04254_),
    .B(_04258_),
    .Y(_04360_));
 sky130_fd_sc_hd__nand2b_1 _09859_ (.A_N(_04259_),
    .B(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__a21o_1 _09860_ (.A1(_04359_),
    .A2(_04360_),
    .B1(_04259_),
    .X(_04362_));
 sky130_fd_sc_hd__nand2_1 _09861_ (.A(_04249_),
    .B(_04252_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand2b_1 _09862_ (.A_N(_04253_),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__a21o_1 _09863_ (.A1(_04362_),
    .A2(_04363_),
    .B1(_04253_),
    .X(_04365_));
 sky130_fd_sc_hd__nand2_1 _09864_ (.A(_04243_),
    .B(_04247_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand2b_1 _09865_ (.A_N(_04248_),
    .B(_04366_),
    .Y(_04368_));
 sky130_fd_sc_hd__a21o_1 _09866_ (.A1(_04365_),
    .A2(_04366_),
    .B1(_04248_),
    .X(_04369_));
 sky130_fd_sc_hd__nand2_1 _09867_ (.A(_04238_),
    .B(_04241_),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2b_1 _09868_ (.A_N(_04242_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__a21o_1 _09869_ (.A1(_04369_),
    .A2(_04370_),
    .B1(_04242_),
    .X(_04372_));
 sky130_fd_sc_hd__nand2_1 _09870_ (.A(_04232_),
    .B(_04236_),
    .Y(_04373_));
 sky130_fd_sc_hd__nand2b_1 _09871_ (.A_N(_04237_),
    .B(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__a21o_1 _09872_ (.A1(_04372_),
    .A2(_04373_),
    .B1(_04237_),
    .X(_04375_));
 sky130_fd_sc_hd__nand2_1 _09873_ (.A(_04227_),
    .B(_04230_),
    .Y(_04376_));
 sky130_fd_sc_hd__nand2b_1 _09874_ (.A_N(_04231_),
    .B(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__a21o_1 _09875_ (.A1(_04375_),
    .A2(_04376_),
    .B1(_04231_),
    .X(_04379_));
 sky130_fd_sc_hd__nand2_1 _09876_ (.A(_04221_),
    .B(_04225_),
    .Y(_04380_));
 sky130_fd_sc_hd__nand2b_1 _09877_ (.A_N(_04226_),
    .B(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__a21o_1 _09878_ (.A1(_04379_),
    .A2(_04380_),
    .B1(_04226_),
    .X(_04382_));
 sky130_fd_sc_hd__nand2_1 _09879_ (.A(_04216_),
    .B(_04219_),
    .Y(_04383_));
 sky130_fd_sc_hd__nand2b_1 _09880_ (.A_N(_04220_),
    .B(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__a21o_1 _09881_ (.A1(_04382_),
    .A2(_04383_),
    .B1(_04220_),
    .X(_04385_));
 sky130_fd_sc_hd__nand2_1 _09882_ (.A(_04210_),
    .B(_04214_),
    .Y(_04386_));
 sky130_fd_sc_hd__nand2b_1 _09883_ (.A_N(_04215_),
    .B(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__a21o_1 _09884_ (.A1(_04385_),
    .A2(_04386_),
    .B1(_04215_),
    .X(_04388_));
 sky130_fd_sc_hd__nand2_1 _09885_ (.A(_04205_),
    .B(_04208_),
    .Y(_04390_));
 sky130_fd_sc_hd__nand2b_1 _09886_ (.A_N(_04209_),
    .B(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__a21o_1 _09887_ (.A1(_04388_),
    .A2(_04390_),
    .B1(_04209_),
    .X(_04392_));
 sky130_fd_sc_hd__nand2_1 _09888_ (.A(_04199_),
    .B(_04203_),
    .Y(_04393_));
 sky130_fd_sc_hd__nand2b_1 _09889_ (.A_N(_04204_),
    .B(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hd__a21o_1 _09890_ (.A1(_04392_),
    .A2(_04393_),
    .B1(_04204_),
    .X(_04395_));
 sky130_fd_sc_hd__nand2_1 _09891_ (.A(_04194_),
    .B(_04197_),
    .Y(_04396_));
 sky130_fd_sc_hd__nand2b_1 _09892_ (.A_N(_04198_),
    .B(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__a21o_1 _09893_ (.A1(_04395_),
    .A2(_04396_),
    .B1(_04198_),
    .X(_04398_));
 sky130_fd_sc_hd__nand2_1 _09894_ (.A(_04188_),
    .B(_04192_),
    .Y(_04399_));
 sky130_fd_sc_hd__nand2b_1 _09895_ (.A_N(_04193_),
    .B(_04399_),
    .Y(_04401_));
 sky130_fd_sc_hd__a21o_1 _09896_ (.A1(_04398_),
    .A2(_04399_),
    .B1(_04193_),
    .X(_04402_));
 sky130_fd_sc_hd__nand2_1 _09897_ (.A(_04183_),
    .B(_04186_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand2b_1 _09898_ (.A_N(_04187_),
    .B(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__a21o_1 _09899_ (.A1(_04402_),
    .A2(_04403_),
    .B1(_04187_),
    .X(_04405_));
 sky130_fd_sc_hd__nand2_1 _09900_ (.A(_04177_),
    .B(_04181_),
    .Y(_04406_));
 sky130_fd_sc_hd__nand2b_1 _09901_ (.A_N(_04182_),
    .B(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__a21o_1 _09902_ (.A1(_04405_),
    .A2(_04406_),
    .B1(_04182_),
    .X(_04408_));
 sky130_fd_sc_hd__nand2_1 _09903_ (.A(_04172_),
    .B(_04175_),
    .Y(_04409_));
 sky130_fd_sc_hd__nand2b_1 _09904_ (.A_N(_04176_),
    .B(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__a21o_1 _09905_ (.A1(_04408_),
    .A2(_04409_),
    .B1(_04176_),
    .X(_04412_));
 sky130_fd_sc_hd__nand2_1 _09906_ (.A(_04134_),
    .B(_04170_),
    .Y(_04413_));
 sky130_fd_sc_hd__nand2b_1 _09907_ (.A_N(_04171_),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__a21o_1 _09908_ (.A1(_04412_),
    .A2(_04413_),
    .B1(_04171_),
    .X(_04415_));
 sky130_fd_sc_hd__nand2_1 _09909_ (.A(net56),
    .B(net25),
    .Y(_04416_));
 sky130_fd_sc_hd__and2b_1 _09910_ (.A_N(_04127_),
    .B(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__and3_1 _09911_ (.A(net56),
    .B(net25),
    .C(_04127_),
    .X(_04418_));
 sky130_fd_sc_hd__or2_1 _09912_ (.A(_04417_),
    .B(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__o211a_1 _09913_ (.A1(_04124_),
    .A2(_04133_),
    .B1(_04419_),
    .C1(_04132_),
    .X(_04420_));
 sky130_fd_sc_hd__or2_1 _09914_ (.A(net24),
    .B(_04167_),
    .X(_04421_));
 sky130_fd_sc_hd__nand2_1 _09915_ (.A(net57),
    .B(_04421_),
    .Y(_04423_));
 sky130_fd_sc_hd__a21oi_1 _09916_ (.A1(net24),
    .A2(_04167_),
    .B1(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__inv_2 _09917_ (.A(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__xnor2_1 _09918_ (.A(_04420_),
    .B(_04424_),
    .Y(_04426_));
 sky130_fd_sc_hd__nand2_1 _09919_ (.A(net25),
    .B(net57),
    .Y(_04427_));
 sky130_fd_sc_hd__o22a_1 _09920_ (.A1(net25),
    .A2(_04423_),
    .B1(_04427_),
    .B2(_04421_),
    .X(_04428_));
 sky130_fd_sc_hd__o22ai_1 _09921_ (.A1(_04420_),
    .A2(_04425_),
    .B1(_04428_),
    .B2(_04417_),
    .Y(_04429_));
 sky130_fd_sc_hd__a21oi_1 _09922_ (.A1(_04415_),
    .A2(_04426_),
    .B1(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__xnor2_1 _09923_ (.A(_02098_),
    .B(_02739_),
    .Y(_04431_));
 sky130_fd_sc_hd__xnor2_1 _09924_ (.A(_01851_),
    .B(_02631_),
    .Y(_04432_));
 sky130_fd_sc_hd__xnor2_1 _09925_ (.A(_01905_),
    .B(_04432_),
    .Y(_04434_));
 sky130_fd_sc_hd__xnor2_1 _09926_ (.A(_02028_),
    .B(_02853_),
    .Y(_04435_));
 sky130_fd_sc_hd__xnor2_1 _09927_ (.A(_04434_),
    .B(_04435_),
    .Y(_04436_));
 sky130_fd_sc_hd__nand2_1 _09928_ (.A(_01760_),
    .B(_01801_),
    .Y(_04437_));
 sky130_fd_sc_hd__o22a_1 _09929_ (.A1(net64),
    .A2(_01848_),
    .B1(_01902_),
    .B2(net63),
    .X(_04438_));
 sky130_fd_sc_hd__o22a_1 _09930_ (.A1(net39),
    .A2(_02026_),
    .B1(_02339_),
    .B2(net35),
    .X(_04439_));
 sky130_fd_sc_hd__xnor2_1 _09931_ (.A(_04438_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__o22a_1 _09932_ (.A1(net41),
    .A2(_02430_),
    .B1(_02528_),
    .B2(net40),
    .X(_04441_));
 sky130_fd_sc_hd__xnor2_1 _09933_ (.A(_02253_),
    .B(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__o22a_1 _09934_ (.A1(net37),
    .A2(_02096_),
    .B1(_02173_),
    .B2(net36),
    .X(_04443_));
 sky130_fd_sc_hd__o22a_1 _09935_ (.A1(net34),
    .A2(_01801_),
    .B1(_01962_),
    .B2(net62),
    .X(_04445_));
 sky130_fd_sc_hd__xor2_1 _09936_ (.A(_04443_),
    .B(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__xnor2_1 _09937_ (.A(_04442_),
    .B(_04446_),
    .Y(_04447_));
 sky130_fd_sc_hd__xnor2_1 _09938_ (.A(_04440_),
    .B(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__xnor2_1 _09939_ (.A(_04437_),
    .B(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__xnor2_1 _09940_ (.A(_01964_),
    .B(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__xnor2_1 _09941_ (.A(_04431_),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__xnor2_1 _09942_ (.A(_03228_),
    .B(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__xnor2_1 _09943_ (.A(_02433_),
    .B(_04436_),
    .Y(_04453_));
 sky130_fd_sc_hd__xnor2_1 _09944_ (.A(_04452_),
    .B(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__and2b_1 _09945_ (.A_N(net42),
    .B(_02530_),
    .X(_04456_));
 sky130_fd_sc_hd__a31o_1 _09946_ (.A1(net42),
    .A2(net25),
    .A3(_02532_),
    .B1(_04456_),
    .X(_04457_));
 sky130_fd_sc_hd__xnor2_1 _09947_ (.A(_04454_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__xor2_1 _09948_ (.A(_02341_),
    .B(_03363_),
    .X(_04459_));
 sky130_fd_sc_hd__nand2_1 _09949_ (.A(_02175_),
    .B(_02255_),
    .Y(_04460_));
 sky130_fd_sc_hd__o21a_1 _09950_ (.A1(net38),
    .A2(_02175_),
    .B1(_04460_),
    .X(_04461_));
 sky130_fd_sc_hd__o22a_1 _09951_ (.A1(net47),
    .A2(_02973_),
    .B1(_03097_),
    .B2(net46),
    .X(_04462_));
 sky130_fd_sc_hd__o22a_1 _09952_ (.A1(net51),
    .A2(_03504_),
    .B1(_03651_),
    .B2(net50),
    .X(_04463_));
 sky130_fd_sc_hd__xor2_1 _09953_ (.A(_04462_),
    .B(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__xnor2_1 _09954_ (.A(_04461_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__xnor2_1 _09955_ (.A(_04459_),
    .B(_04465_),
    .Y(_04467_));
 sky130_fd_sc_hd__xnor2_1 _09956_ (.A(_04458_),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__nor2_1 _09957_ (.A(net45),
    .B(_02742_),
    .Y(_04469_));
 sky130_fd_sc_hd__a31o_1 _09958_ (.A1(net45),
    .A2(net25),
    .A3(_02743_),
    .B1(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__o22a_1 _09959_ (.A1(net53),
    .A2(_03803_),
    .B1(_03963_),
    .B2(net52),
    .X(_04471_));
 sky130_fd_sc_hd__xnor2_1 _09960_ (.A(_04126_),
    .B(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__xnor2_1 _09961_ (.A(_04470_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__xnor2_1 _09962_ (.A(_04468_),
    .B(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__xnor2_1 _09963_ (.A(_03365_),
    .B(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__xnor2_1 _09964_ (.A(_02975_),
    .B(_04416_),
    .Y(_04476_));
 sky130_fd_sc_hd__nand2_1 _09965_ (.A(_03099_),
    .B(_03230_),
    .Y(_04478_));
 sky130_fd_sc_hd__o21a_1 _09966_ (.A1(net48),
    .A2(_03099_),
    .B1(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__xnor2_1 _09967_ (.A(_04476_),
    .B(_04479_),
    .Y(_04480_));
 sky130_fd_sc_hd__xnor2_1 _09968_ (.A(_04475_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__nand2_1 _09969_ (.A(_03506_),
    .B(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__o221a_1 _09970_ (.A1(net25),
    .A2(_04423_),
    .B1(_04481_),
    .B2(_03506_),
    .C1(_04482_),
    .X(_04483_));
 sky130_fd_sc_hd__and2b_1 _09971_ (.A_N(net52),
    .B(_03654_),
    .X(_04484_));
 sky130_fd_sc_hd__a31o_1 _09972_ (.A1(net52),
    .A2(net25),
    .A3(_03655_),
    .B1(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__nand2_1 _09973_ (.A(_03965_),
    .B(_04128_),
    .Y(_04486_));
 sky130_fd_sc_hd__o21ai_1 _09974_ (.A1(net54),
    .A2(_03965_),
    .B1(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__xnor2_1 _09975_ (.A(_04485_),
    .B(_04487_),
    .Y(_04489_));
 sky130_fd_sc_hd__xnor2_1 _09976_ (.A(_04483_),
    .B(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__xnor2_1 _09977_ (.A(_04418_),
    .B(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__xnor2_1 _09978_ (.A(_04430_),
    .B(_04491_),
    .Y(\genblk2[30].rca1.ripple_adders[31].fa.sum ));
 sky130_fd_sc_hd__a21boi_1 _09979_ (.A1(_04417_),
    .A2(_04428_),
    .B1_N(_04430_),
    .Y(\genblk2[30].rca1.ripple_adders[30].fa.sum ));
 sky130_fd_sc_hd__xor2_1 _09980_ (.A(_04415_),
    .B(_04426_),
    .X(\genblk2[30].rca1.ripple_adders[29].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09981_ (.A(_04412_),
    .B(_04414_),
    .Y(\genblk2[30].rca1.ripple_adders[28].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09982_ (.A(_04408_),
    .B(_04410_),
    .Y(\genblk2[30].rca1.ripple_adders[27].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09983_ (.A(_04405_),
    .B(_04407_),
    .Y(\genblk2[30].rca1.ripple_adders[26].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09984_ (.A(_04402_),
    .B(_04404_),
    .Y(\genblk2[30].rca1.ripple_adders[25].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09985_ (.A(_04398_),
    .B(_04401_),
    .Y(\genblk2[30].rca1.ripple_adders[24].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09986_ (.A(_04395_),
    .B(_04397_),
    .Y(\genblk2[30].rca1.ripple_adders[23].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09987_ (.A(_04392_),
    .B(_04394_),
    .Y(\genblk2[30].rca1.ripple_adders[22].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09988_ (.A(_04388_),
    .B(_04391_),
    .Y(\genblk2[30].rca1.ripple_adders[21].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09989_ (.A(_04385_),
    .B(_04387_),
    .Y(\genblk2[30].rca1.ripple_adders[20].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09990_ (.A(_04382_),
    .B(_04384_),
    .Y(\genblk2[30].rca1.ripple_adders[19].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09991_ (.A(_04379_),
    .B(_04381_),
    .Y(\genblk2[30].rca1.ripple_adders[18].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09992_ (.A(_04375_),
    .B(_04377_),
    .Y(\genblk2[30].rca1.ripple_adders[17].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09993_ (.A(_04372_),
    .B(_04374_),
    .Y(\genblk2[30].rca1.ripple_adders[16].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09994_ (.A(_04369_),
    .B(_04371_),
    .Y(\genblk2[30].rca1.ripple_adders[15].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09995_ (.A(_04365_),
    .B(_04368_),
    .Y(\genblk2[30].rca1.ripple_adders[14].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09996_ (.A(_04362_),
    .B(_04364_),
    .Y(\genblk2[30].rca1.ripple_adders[13].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09997_ (.A(_04359_),
    .B(_04361_),
    .Y(\genblk2[30].rca1.ripple_adders[12].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09998_ (.A(_04355_),
    .B(_04358_),
    .Y(\genblk2[30].rca1.ripple_adders[11].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _09999_ (.A(_04352_),
    .B(_04354_),
    .Y(\genblk2[30].rca1.ripple_adders[10].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _10000_ (.A(_04349_),
    .B(_04351_),
    .Y(\genblk2[30].rca1.ripple_adders[9].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _10001_ (.A(_04346_),
    .B(_04348_),
    .Y(\genblk2[30].rca1.ripple_adders[8].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _10002_ (.A(_04342_),
    .B(_04344_),
    .Y(\genblk2[30].rca1.ripple_adders[7].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _10003_ (.A(_04339_),
    .B(_04341_),
    .Y(\genblk2[30].rca1.ripple_adders[6].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _10004_ (.A(_04336_),
    .B(_04338_),
    .Y(\genblk2[30].rca1.ripple_adders[5].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _10005_ (.A(_04332_),
    .B(_04335_),
    .Y(\genblk2[30].rca1.ripple_adders[4].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _10006_ (.A(_04329_),
    .B(_04331_),
    .Y(\genblk2[30].rca1.ripple_adders[3].fa.sum ));
 sky130_fd_sc_hd__xnor2_1 _10007_ (.A(_04326_),
    .B(_04328_),
    .Y(\genblk2[30].rca1.ripple_adders[2].fa.sum ));
 sky130_fd_sc_hd__xor2_1 _10008_ (.A(_04324_),
    .B(_04325_),
    .X(\genblk2[30].rca1.ripple_adders[1].fa.sum ));
 sky130_fd_sc_hd__xor2_1 _10009_ (.A(_01634_),
    .B(_04322_),
    .X(\genblk2[30].rca1.ripple_adders[0].fa.sum ));
 sky130_fd_sc_hd__a22o_1 _10010_ (.A1(net12),
    .A2(net33),
    .B1(net44),
    .B2(net1),
    .X(_04495_));
 sky130_fd_sc_hd__o21a_1 _10011_ (.A1(_00384_),
    .A2(_00395_),
    .B1(_04495_),
    .X(\genblk2[10].rca.ripple_adders[1].fa.a ));
 sky130_fd_sc_hd__and3_1 _10012_ (.A(_00287_),
    .B(_00329_),
    .C(_00340_),
    .X(_04496_));
 sky130_fd_sc_hd__nor2_1 _10013_ (.A(_00351_),
    .B(_04496_),
    .Y(\genblk2[10].rca.ripple_adders[2].fa.a ));
 sky130_fd_sc_hd__a21oi_1 _10014_ (.A1(net1),
    .A2(net58),
    .B1(_00471_),
    .Y(_04497_));
 sky130_fd_sc_hd__nor2_1 _10015_ (.A(_00482_),
    .B(_04497_),
    .Y(\genblk2[10].rca.ripple_adders[3].fa.a ));
 sky130_fd_sc_hd__a21oi_1 _10016_ (.A1(net1),
    .A2(net59),
    .B1(_00635_),
    .Y(_04499_));
 sky130_fd_sc_hd__nor2_1 _10017_ (.A(_00646_),
    .B(_04499_),
    .Y(\genblk2[10].rca.ripple_adders[4].fa.a ));
 sky130_fd_sc_hd__a21oi_1 _10018_ (.A1(net1),
    .A2(net60),
    .B1(_00864_),
    .Y(_04500_));
 sky130_fd_sc_hd__nor2_1 _10019_ (.A(_00875_),
    .B(_04500_),
    .Y(\genblk2[10].rca.ripple_adders[5].fa.a ));
 sky130_fd_sc_hd__a21oi_1 _10020_ (.A1(net1),
    .A2(net61),
    .B1(_01149_),
    .Y(_04501_));
 sky130_fd_sc_hd__nor2_1 _10021_ (.A(_01159_),
    .B(_04501_),
    .Y(\genblk2[10].rca.ripple_adders[6].fa.a ));
 sky130_fd_sc_hd__a21oi_1 _10022_ (.A1(net1),
    .A2(net62),
    .B1(_01487_),
    .Y(_04502_));
 sky130_fd_sc_hd__nor2_1 _10023_ (.A(_01498_),
    .B(_04502_),
    .Y(\genblk2[10].rca.ripple_adders[7].fa.a ));
 sky130_fd_sc_hd__a21oi_1 _10024_ (.A1(net1),
    .A2(net63),
    .B1(_01882_),
    .Y(_04503_));
 sky130_fd_sc_hd__nor2_1 _10025_ (.A(_01893_),
    .B(_04503_),
    .Y(\genblk2[10].rca.ripple_adders[8].fa.a ));
 sky130_fd_sc_hd__a21oi_1 _10026_ (.A1(net64),
    .A2(net1),
    .B1(_02333_),
    .Y(_04505_));
 sky130_fd_sc_hd__nor2_1 _10027_ (.A(_02344_),
    .B(_04505_),
    .Y(\genblk2[10].rca.ripple_adders[9].fa.a ));
 sky130_fd_sc_hd__a21oi_1 _10028_ (.A1(net34),
    .A2(net1),
    .B1(_02839_),
    .Y(_04506_));
 sky130_fd_sc_hd__nor2_1 _10029_ (.A(_02850_),
    .B(_04506_),
    .Y(\genblk2[10].rca.ripple_adders[10].fa.a ));
 sky130_fd_sc_hd__a21oi_1 _10030_ (.A1(net35),
    .A2(net1),
    .B1(_03400_),
    .Y(_04507_));
 sky130_fd_sc_hd__nor2_1 _10031_ (.A(_03411_),
    .B(_04507_),
    .Y(\genblk2[10].rca.ripple_adders[11].fa.sum ));
 sky130_fd_sc_hd__buf_1 _10032_ (.A(\genblk2[10].rca.ripple_adders[0].fa.a ),
    .X(net65));
 sky130_fd_sc_hd__buf_1 _10033_ (.A(\genblk2[10].rca.ripple_adders[1].fa.a ),
    .X(net76));
 sky130_fd_sc_hd__buf_1 _10034_ (.A(\genblk2[10].rca.ripple_adders[2].fa.a ),
    .X(net87));
 sky130_fd_sc_hd__buf_1 _10035_ (.A(\genblk2[10].rca.ripple_adders[3].fa.a ),
    .X(net98));
 sky130_fd_sc_hd__buf_1 _10036_ (.A(\genblk2[10].rca.ripple_adders[4].fa.a ),
    .X(net109));
 sky130_fd_sc_hd__buf_1 _10037_ (.A(\genblk2[10].rca.ripple_adders[5].fa.a ),
    .X(net120));
 sky130_fd_sc_hd__buf_1 _10038_ (.A(\genblk2[10].rca.ripple_adders[6].fa.a ),
    .X(net125));
 sky130_fd_sc_hd__buf_1 _10039_ (.A(\genblk2[10].rca.ripple_adders[7].fa.a ),
    .X(net126));
 sky130_fd_sc_hd__buf_1 _10040_ (.A(\genblk2[10].rca.ripple_adders[8].fa.a ),
    .X(net127));
 sky130_fd_sc_hd__buf_1 _10041_ (.A(\genblk2[10].rca.ripple_adders[9].fa.a ),
    .X(net128));
 sky130_fd_sc_hd__buf_1 _10042_ (.A(\genblk2[10].rca.ripple_adders[10].fa.a ),
    .X(net66));
 sky130_fd_sc_hd__buf_1 _10043_ (.A(\genblk2[10].rca.ripple_adders[11].fa.sum ),
    .X(net67));
 sky130_fd_sc_hd__buf_1 _10044_ (.A(\genblk2[11].rca.ripple_adders[12].fa.sum ),
    .X(net68));
 sky130_fd_sc_hd__buf_1 _10045_ (.A(\genblk2[12].rca.ripple_adders[13].fa.sum ),
    .X(net69));
 sky130_fd_sc_hd__buf_1 _10046_ (.A(\genblk2[13].rca.ripple_adders[14].fa.sum ),
    .X(net70));
 sky130_fd_sc_hd__buf_1 _10047_ (.A(\genblk2[14].rca.ripple_adders[15].fa.sum ),
    .X(net71));
 sky130_fd_sc_hd__buf_1 _10048_ (.A(\genblk2[15].rca.ripple_adders[16].fa.sum ),
    .X(net72));
 sky130_fd_sc_hd__buf_1 _10049_ (.A(\genblk2[16].rca.ripple_adders[17].fa.sum ),
    .X(net73));
 sky130_fd_sc_hd__buf_1 _10050_ (.A(\genblk2[17].rca.ripple_adders[18].fa.sum ),
    .X(net74));
 sky130_fd_sc_hd__buf_1 _10051_ (.A(\genblk2[18].rca.ripple_adders[19].fa.sum ),
    .X(net75));
 sky130_fd_sc_hd__buf_1 _10052_ (.A(\genblk2[19].rca.ripple_adders[20].fa.sum ),
    .X(net77));
 sky130_fd_sc_hd__buf_1 _10053_ (.A(\genblk2[20].rca.ripple_adders[21].fa.sum ),
    .X(net78));
 sky130_fd_sc_hd__buf_1 _10054_ (.A(\genblk2[21].rca.ripple_adders[22].fa.sum ),
    .X(net79));
 sky130_fd_sc_hd__buf_1 _10055_ (.A(\genblk2[22].rca.ripple_adders[23].fa.sum ),
    .X(net80));
 sky130_fd_sc_hd__buf_1 _10056_ (.A(\genblk2[23].rca.ripple_adders[24].fa.sum ),
    .X(net81));
 sky130_fd_sc_hd__buf_1 _10057_ (.A(\genblk2[24].rca.ripple_adders[25].fa.sum ),
    .X(net82));
 sky130_fd_sc_hd__buf_1 _10058_ (.A(\genblk2[25].rca.ripple_adders[26].fa.sum ),
    .X(net83));
 sky130_fd_sc_hd__buf_1 _10059_ (.A(\genblk2[26].rca.ripple_adders[27].fa.sum ),
    .X(net84));
 sky130_fd_sc_hd__buf_1 _10060_ (.A(\genblk2[27].rca.ripple_adders[28].fa.sum ),
    .X(net85));
 sky130_fd_sc_hd__buf_1 _10061_ (.A(\genblk2[28].rca.ripple_adders[29].fa.sum ),
    .X(net86));
 sky130_fd_sc_hd__buf_1 _10062_ (.A(\genblk2[29].rca.ripple_adders[30].fa.sum ),
    .X(net88));
 sky130_fd_sc_hd__buf_1 _10063_ (.A(\genblk2[30].rca.ripple_adders[31].fa.sum ),
    .X(net89));
 sky130_fd_sc_hd__buf_1 _10064_ (.A(\genblk2[30].rca1.ripple_adders[0].fa.sum ),
    .X(net90));
 sky130_fd_sc_hd__buf_1 _10065_ (.A(\genblk2[30].rca1.ripple_adders[1].fa.sum ),
    .X(net91));
 sky130_fd_sc_hd__buf_1 _10066_ (.A(\genblk2[30].rca1.ripple_adders[2].fa.sum ),
    .X(net92));
 sky130_fd_sc_hd__buf_1 _10067_ (.A(\genblk2[30].rca1.ripple_adders[3].fa.sum ),
    .X(net93));
 sky130_fd_sc_hd__buf_1 _10068_ (.A(\genblk2[30].rca1.ripple_adders[4].fa.sum ),
    .X(net94));
 sky130_fd_sc_hd__buf_1 _10069_ (.A(\genblk2[30].rca1.ripple_adders[5].fa.sum ),
    .X(net95));
 sky130_fd_sc_hd__buf_1 _10070_ (.A(\genblk2[30].rca1.ripple_adders[6].fa.sum ),
    .X(net96));
 sky130_fd_sc_hd__buf_1 _10071_ (.A(\genblk2[30].rca1.ripple_adders[7].fa.sum ),
    .X(net97));
 sky130_fd_sc_hd__buf_1 _10072_ (.A(\genblk2[30].rca1.ripple_adders[8].fa.sum ),
    .X(net99));
 sky130_fd_sc_hd__buf_1 _10073_ (.A(\genblk2[30].rca1.ripple_adders[9].fa.sum ),
    .X(net100));
 sky130_fd_sc_hd__buf_1 _10074_ (.A(\genblk2[30].rca1.ripple_adders[10].fa.sum ),
    .X(net101));
 sky130_fd_sc_hd__buf_1 _10075_ (.A(\genblk2[30].rca1.ripple_adders[11].fa.sum ),
    .X(net102));
 sky130_fd_sc_hd__buf_1 _10076_ (.A(\genblk2[30].rca1.ripple_adders[12].fa.sum ),
    .X(net103));
 sky130_fd_sc_hd__buf_1 _10077_ (.A(\genblk2[30].rca1.ripple_adders[13].fa.sum ),
    .X(net104));
 sky130_fd_sc_hd__buf_1 _10078_ (.A(\genblk2[30].rca1.ripple_adders[14].fa.sum ),
    .X(net105));
 sky130_fd_sc_hd__buf_1 _10079_ (.A(\genblk2[30].rca1.ripple_adders[15].fa.sum ),
    .X(net106));
 sky130_fd_sc_hd__buf_1 _10080_ (.A(\genblk2[30].rca1.ripple_adders[16].fa.sum ),
    .X(net107));
 sky130_fd_sc_hd__buf_1 _10081_ (.A(\genblk2[30].rca1.ripple_adders[17].fa.sum ),
    .X(net108));
 sky130_fd_sc_hd__buf_1 _10082_ (.A(\genblk2[30].rca1.ripple_adders[18].fa.sum ),
    .X(net110));
 sky130_fd_sc_hd__buf_1 _10083_ (.A(\genblk2[30].rca1.ripple_adders[19].fa.sum ),
    .X(net111));
 sky130_fd_sc_hd__buf_1 _10084_ (.A(\genblk2[30].rca1.ripple_adders[20].fa.sum ),
    .X(net112));
 sky130_fd_sc_hd__buf_1 _10085_ (.A(\genblk2[30].rca1.ripple_adders[21].fa.sum ),
    .X(net113));
 sky130_fd_sc_hd__buf_1 _10086_ (.A(\genblk2[30].rca1.ripple_adders[22].fa.sum ),
    .X(net114));
 sky130_fd_sc_hd__buf_1 _10087_ (.A(\genblk2[30].rca1.ripple_adders[23].fa.sum ),
    .X(net115));
 sky130_fd_sc_hd__buf_1 _10088_ (.A(\genblk2[30].rca1.ripple_adders[24].fa.sum ),
    .X(net116));
 sky130_fd_sc_hd__buf_1 _10089_ (.A(\genblk2[30].rca1.ripple_adders[25].fa.sum ),
    .X(net117));
 sky130_fd_sc_hd__buf_1 _10090_ (.A(\genblk2[30].rca1.ripple_adders[26].fa.sum ),
    .X(net118));
 sky130_fd_sc_hd__buf_1 _10091_ (.A(\genblk2[30].rca1.ripple_adders[27].fa.sum ),
    .X(net119));
 sky130_fd_sc_hd__buf_1 _10092_ (.A(\genblk2[30].rca1.ripple_adders[28].fa.sum ),
    .X(net121));
 sky130_fd_sc_hd__buf_1 _10093_ (.A(\genblk2[30].rca1.ripple_adders[29].fa.sum ),
    .X(net122));
 sky130_fd_sc_hd__buf_1 _10094_ (.A(\genblk2[30].rca1.ripple_adders[30].fa.sum ),
    .X(net123));
 sky130_fd_sc_hd__buf_1 _10095_ (.A(\genblk2[30].rca1.ripple_adders[31].fa.sum ),
    .X(net124));
 sky130_fd_sc_hd__buf_12 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_16 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_16 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_16 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_16 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_16 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_16 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_16 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_16 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_16 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_16 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_16 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_16 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_16 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_12 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_12 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_16 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_16 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_16 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_16 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_16 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_16 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_16 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_12 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_16 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_16 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_16 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_16 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_16 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_16 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_16 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_16 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_12 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_16 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_16 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_16 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_8 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_8 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_8 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_8 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_8 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_16 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_8 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_12 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_16 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_8 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_8 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_16 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_8 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_8 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_16 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_12 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_16 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_16 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_12 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_16 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_6 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_12 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_12 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_12 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_12 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_12 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_12 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_16 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_16 output65 (.A(net65),
    .X(z[0]));
 sky130_fd_sc_hd__clkbuf_16 output66 (.A(net66),
    .X(z[10]));
 sky130_fd_sc_hd__clkbuf_16 output67 (.A(net67),
    .X(z[11]));
 sky130_fd_sc_hd__clkbuf_16 output68 (.A(net68),
    .X(z[12]));
 sky130_fd_sc_hd__clkbuf_16 output69 (.A(net69),
    .X(z[13]));
 sky130_fd_sc_hd__clkbuf_16 output70 (.A(net70),
    .X(z[14]));
 sky130_fd_sc_hd__clkbuf_16 output71 (.A(net71),
    .X(z[15]));
 sky130_fd_sc_hd__clkbuf_16 output72 (.A(net72),
    .X(z[16]));
 sky130_fd_sc_hd__clkbuf_16 output73 (.A(net73),
    .X(z[17]));
 sky130_fd_sc_hd__clkbuf_16 output74 (.A(net74),
    .X(z[18]));
 sky130_fd_sc_hd__clkbuf_16 output75 (.A(net75),
    .X(z[19]));
 sky130_fd_sc_hd__clkbuf_16 output76 (.A(net76),
    .X(z[1]));
 sky130_fd_sc_hd__clkbuf_16 output77 (.A(net77),
    .X(z[20]));
 sky130_fd_sc_hd__clkbuf_16 output78 (.A(net78),
    .X(z[21]));
 sky130_fd_sc_hd__clkbuf_16 output79 (.A(net79),
    .X(z[22]));
 sky130_fd_sc_hd__clkbuf_16 output80 (.A(net80),
    .X(z[23]));
 sky130_fd_sc_hd__clkbuf_16 output81 (.A(net81),
    .X(z[24]));
 sky130_fd_sc_hd__clkbuf_16 output82 (.A(net82),
    .X(z[25]));
 sky130_fd_sc_hd__clkbuf_16 output83 (.A(net83),
    .X(z[26]));
 sky130_fd_sc_hd__clkbuf_16 output84 (.A(net84),
    .X(z[27]));
 sky130_fd_sc_hd__clkbuf_16 output85 (.A(net85),
    .X(z[28]));
 sky130_fd_sc_hd__clkbuf_16 output86 (.A(net86),
    .X(z[29]));
 sky130_fd_sc_hd__clkbuf_16 output87 (.A(net87),
    .X(z[2]));
 sky130_fd_sc_hd__clkbuf_16 output88 (.A(net88),
    .X(z[30]));
 sky130_fd_sc_hd__clkbuf_16 output89 (.A(net89),
    .X(z[31]));
 sky130_fd_sc_hd__clkbuf_16 output90 (.A(net90),
    .X(z[32]));
 sky130_fd_sc_hd__clkbuf_16 output91 (.A(net91),
    .X(z[33]));
 sky130_fd_sc_hd__clkbuf_16 output92 (.A(net92),
    .X(z[34]));
 sky130_fd_sc_hd__clkbuf_16 output93 (.A(net93),
    .X(z[35]));
 sky130_fd_sc_hd__clkbuf_16 output94 (.A(net94),
    .X(z[36]));
 sky130_fd_sc_hd__clkbuf_16 output95 (.A(net95),
    .X(z[37]));
 sky130_fd_sc_hd__clkbuf_16 output96 (.A(net96),
    .X(z[38]));
 sky130_fd_sc_hd__clkbuf_16 output97 (.A(net97),
    .X(z[39]));
 sky130_fd_sc_hd__clkbuf_16 output98 (.A(net98),
    .X(z[3]));
 sky130_fd_sc_hd__clkbuf_16 output99 (.A(net99),
    .X(z[40]));
 sky130_fd_sc_hd__clkbuf_16 output100 (.A(net100),
    .X(z[41]));
 sky130_fd_sc_hd__clkbuf_16 output101 (.A(net101),
    .X(z[42]));
 sky130_fd_sc_hd__clkbuf_16 output102 (.A(net102),
    .X(z[43]));
 sky130_fd_sc_hd__clkbuf_16 output103 (.A(net103),
    .X(z[44]));
 sky130_fd_sc_hd__clkbuf_16 output104 (.A(net104),
    .X(z[45]));
 sky130_fd_sc_hd__clkbuf_16 output105 (.A(net105),
    .X(z[46]));
 sky130_fd_sc_hd__clkbuf_16 output106 (.A(net106),
    .X(z[47]));
 sky130_fd_sc_hd__clkbuf_16 output107 (.A(net107),
    .X(z[48]));
 sky130_fd_sc_hd__clkbuf_16 output108 (.A(net108),
    .X(z[49]));
 sky130_fd_sc_hd__clkbuf_16 output109 (.A(net109),
    .X(z[4]));
 sky130_fd_sc_hd__clkbuf_16 output110 (.A(net110),
    .X(z[50]));
 sky130_fd_sc_hd__clkbuf_16 output111 (.A(net111),
    .X(z[51]));
 sky130_fd_sc_hd__clkbuf_16 output112 (.A(net112),
    .X(z[52]));
 sky130_fd_sc_hd__clkbuf_16 output113 (.A(net113),
    .X(z[53]));
 sky130_fd_sc_hd__clkbuf_16 output114 (.A(net114),
    .X(z[54]));
 sky130_fd_sc_hd__clkbuf_16 output115 (.A(net115),
    .X(z[55]));
 sky130_fd_sc_hd__clkbuf_16 output116 (.A(net116),
    .X(z[56]));
 sky130_fd_sc_hd__clkbuf_16 output117 (.A(net117),
    .X(z[57]));
 sky130_fd_sc_hd__clkbuf_16 output118 (.A(net118),
    .X(z[58]));
 sky130_fd_sc_hd__clkbuf_16 output119 (.A(net119),
    .X(z[59]));
 sky130_fd_sc_hd__clkbuf_16 output120 (.A(net120),
    .X(z[5]));
 sky130_fd_sc_hd__clkbuf_16 output121 (.A(net121),
    .X(z[60]));
 sky130_fd_sc_hd__clkbuf_16 output122 (.A(net122),
    .X(z[61]));
 sky130_fd_sc_hd__clkbuf_16 output123 (.A(net123),
    .X(z[62]));
 sky130_fd_sc_hd__clkbuf_16 output124 (.A(net124),
    .X(z[63]));
 sky130_fd_sc_hd__clkbuf_16 output125 (.A(net125),
    .X(z[6]));
 sky130_fd_sc_hd__clkbuf_16 output126 (.A(net126),
    .X(z[7]));
 sky130_fd_sc_hd__clkbuf_16 output127 (.A(net127),
    .X(z[8]));
 sky130_fd_sc_hd__clkbuf_16 output128 (.A(net128),
    .X(z[9]));
endmodule
