module FP_ALU_route (sel,
    in1,
    in2,
    result);
 input sel;
 input [31:0] in1;
 input [31:0] in2;
 output [31:0] result;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 sky130_fd_sc_hd__clkinv_4 _4209_ (.A(net27),
    .Y(_4187_));
 sky130_fd_sc_hd__clkinv_4 _4210_ (.A(net1),
    .Y(_4198_));
 sky130_fd_sc_hd__inv_2 _4211_ (.A(net13),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _4212_ (.A(net3),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _4213_ (.A(net58),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _4214_ (.A(net60),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _4215_ (.A(net64),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _4216_ (.A(net35),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _4217_ (.A(net36),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _4218_ (.A(net37),
    .Y(_0077_));
 sky130_fd_sc_hd__clkinv_4 _4219_ (.A(net39),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _4220_ (.A(net40),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _4221_ (.A(net47),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _4222_ (.A(net16),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _4223_ (.A(net18),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _4224_ (.A(net22),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _4225_ (.A(net48),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _4226_ (.A(net51),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _4227_ (.A(net65),
    .Y(_0176_));
 sky130_fd_sc_hd__and4_1 _4228_ (.A(net51),
    .B(net54),
    .C(net53),
    .D(net56),
    .X(_0187_));
 sky130_fd_sc_hd__and4_1 _4229_ (.A(net48),
    .B(net50),
    .C(net49),
    .D(net52),
    .X(_0198_));
 sky130_fd_sc_hd__nand2_1 _4230_ (.A(_0187_),
    .B(_0198_),
    .Y(_0209_));
 sky130_fd_sc_hd__or4_2 _4231_ (.A(net59),
    .B(net60),
    .C(net61),
    .D(net62),
    .X(_0220_));
 sky130_fd_sc_hd__or4_1 _4232_ (.A(net44),
    .B(net33),
    .C(net55),
    .D(net58),
    .X(_0231_));
 sky130_fd_sc_hd__or4_1 _4233_ (.A(net36),
    .B(net37),
    .C(net38),
    .D(net39),
    .X(_0242_));
 sky130_fd_sc_hd__or4_1 _4234_ (.A(net63),
    .B(net64),
    .C(net34),
    .D(net35),
    .X(_0253_));
 sky130_fd_sc_hd__or4_1 _4235_ (.A(net40),
    .B(net41),
    .C(net42),
    .D(net43),
    .X(_0264_));
 sky130_fd_sc_hd__or4_1 _4236_ (.A(net45),
    .B(net46),
    .C(net47),
    .D(_0264_),
    .X(_0275_));
 sky130_fd_sc_hd__or3_2 _4237_ (.A(_0242_),
    .B(_0253_),
    .C(_0275_),
    .X(_0286_));
 sky130_fd_sc_hd__nor3_1 _4238_ (.A(_0220_),
    .B(_0231_),
    .C(_0286_),
    .Y(_0297_));
 sky130_fd_sc_hd__or4_2 _4239_ (.A(_0209_),
    .B(_0220_),
    .C(_0231_),
    .D(_0286_),
    .X(_0308_));
 sky130_fd_sc_hd__or4_1 _4240_ (.A(net12),
    .B(net1),
    .C(net15),
    .D(net14),
    .X(_0319_));
 sky130_fd_sc_hd__or4_1 _4241_ (.A(net28),
    .B(net27),
    .C(net26),
    .D(net23),
    .X(_0330_));
 sky130_fd_sc_hd__or4_1 _4242_ (.A(net8),
    .B(net7),
    .C(net6),
    .D(net5),
    .X(_0341_));
 sky130_fd_sc_hd__or4_1 _4243_ (.A(net13),
    .B(net11),
    .C(net10),
    .D(_0341_),
    .X(_0352_));
 sky130_fd_sc_hd__or3_1 _4244_ (.A(net31),
    .B(net30),
    .C(net29),
    .X(_0363_));
 sky130_fd_sc_hd__or4_1 _4245_ (.A(net4),
    .B(net3),
    .C(net2),
    .D(net32),
    .X(_0374_));
 sky130_fd_sc_hd__or4_1 _4246_ (.A(_0319_),
    .B(_0330_),
    .C(_0363_),
    .D(_0374_),
    .X(_0385_));
 sky130_fd_sc_hd__nor3_2 _4247_ (.A(net9),
    .B(_0352_),
    .C(_0385_),
    .Y(_0396_));
 sky130_fd_sc_hd__and4_1 _4248_ (.A(net19),
    .B(net21),
    .C(net22),
    .D(net24),
    .X(_0407_));
 sky130_fd_sc_hd__and4_1 _4249_ (.A(net16),
    .B(net18),
    .C(net17),
    .D(net20),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_1 _4250_ (.A(_0407_),
    .B(_0418_),
    .Y(_0429_));
 sky130_fd_sc_hd__inv_2 _4251_ (.A(_0429_),
    .Y(_0440_));
 sky130_fd_sc_hd__nand2_2 _4252_ (.A(_0396_),
    .B(_0440_),
    .Y(_0451_));
 sky130_fd_sc_hd__nand2_1 _4253_ (.A(_0308_),
    .B(_0451_),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2b_2 _4254_ (.A_N(net56),
    .B(net24),
    .Y(_0473_));
 sky130_fd_sc_hd__inv_2 _4255_ (.A(_0473_),
    .Y(_0484_));
 sky130_fd_sc_hd__and2b_1 _4256_ (.A_N(net24),
    .B(net56),
    .X(_0495_));
 sky130_fd_sc_hd__xor2_2 _4257_ (.A(net22),
    .B(net54),
    .X(_0506_));
 sky130_fd_sc_hd__nand2b_1 _4258_ (.A_N(net53),
    .B(net21),
    .Y(_0517_));
 sky130_fd_sc_hd__and2b_1 _4259_ (.A_N(net21),
    .B(net53),
    .X(_0528_));
 sky130_fd_sc_hd__nand2b_1 _4260_ (.A_N(net21),
    .B(net53),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2b_1 _4261_ (.A_N(net20),
    .B(net52),
    .Y(_0550_));
 sky130_fd_sc_hd__nand2b_1 _4262_ (.A_N(net52),
    .B(net20),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_2 _4263_ (.A(_0550_),
    .B(_0561_),
    .Y(_0572_));
 sky130_fd_sc_hd__nand2b_1 _4264_ (.A_N(net49),
    .B(net17),
    .Y(_0583_));
 sky130_fd_sc_hd__and2b_1 _4265_ (.A_N(net17),
    .B(net49),
    .X(_0594_));
 sky130_fd_sc_hd__nand2b_1 _4266_ (.A_N(net17),
    .B(net49),
    .Y(_0605_));
 sky130_fd_sc_hd__nand2_2 _4267_ (.A(_0583_),
    .B(_0605_),
    .Y(_0616_));
 sky130_fd_sc_hd__a21oi_1 _4268_ (.A1(net16),
    .A2(_0154_),
    .B1(_0616_),
    .Y(_0627_));
 sky130_fd_sc_hd__xnor2_4 _4269_ (.A(net16),
    .B(net48),
    .Y(_0638_));
 sky130_fd_sc_hd__clkinv_4 _4270_ (.A(_0638_),
    .Y(_0649_));
 sky130_fd_sc_hd__nor2_1 _4271_ (.A(_0132_),
    .B(net50),
    .Y(_0660_));
 sky130_fd_sc_hd__and2_1 _4272_ (.A(_0132_),
    .B(net50),
    .X(_0671_));
 sky130_fd_sc_hd__or2_2 _4273_ (.A(_0660_),
    .B(_0671_),
    .X(_0682_));
 sky130_fd_sc_hd__xor2_4 _4274_ (.A(net19),
    .B(net51),
    .X(_0693_));
 sky130_fd_sc_hd__or4_4 _4275_ (.A(_0616_),
    .B(_0649_),
    .C(_0682_),
    .D(_0693_),
    .X(_0704_));
 sky130_fd_sc_hd__a311o_1 _4276_ (.A1(_0121_),
    .A2(net48),
    .A3(_0583_),
    .B1(_0594_),
    .C1(_0671_),
    .X(_0715_));
 sky130_fd_sc_hd__and2b_1 _4277_ (.A_N(_0660_),
    .B(_0715_),
    .X(_0726_));
 sky130_fd_sc_hd__a21bo_1 _4278_ (.A1(net19),
    .A2(_0165_),
    .B1_N(_0726_),
    .X(_0737_));
 sky130_fd_sc_hd__o211a_2 _4279_ (.A1(net19),
    .A2(_0165_),
    .B1(_0704_),
    .C1(_0737_),
    .X(_0748_));
 sky130_fd_sc_hd__o21ai_1 _4280_ (.A1(_0572_),
    .A2(_0748_),
    .B1(_0550_),
    .Y(_0759_));
 sky130_fd_sc_hd__a21o_1 _4281_ (.A1(_0517_),
    .A2(_0759_),
    .B1(_0528_),
    .X(_0770_));
 sky130_fd_sc_hd__and2b_1 _4282_ (.A_N(_0506_),
    .B(_0770_),
    .X(_0781_));
 sky130_fd_sc_hd__a21o_1 _4283_ (.A1(_0143_),
    .A2(net54),
    .B1(_0781_),
    .X(_0792_));
 sky130_fd_sc_hd__a21o_4 _4284_ (.A1(_0473_),
    .A2(_0792_),
    .B1(_0495_),
    .X(_0803_));
 sky130_fd_sc_hd__a21oi_4 _4285_ (.A1(_0473_),
    .A2(_0792_),
    .B1(_0495_),
    .Y(_0814_));
 sky130_fd_sc_hd__nand2_2 _4286_ (.A(_0517_),
    .B(_0539_),
    .Y(_0825_));
 sky130_fd_sc_hd__nor2_1 _4287_ (.A(_0484_),
    .B(_0495_),
    .Y(_0836_));
 sky130_fd_sc_hd__or4b_2 _4288_ (.A(_0506_),
    .B(_0572_),
    .C(_0825_),
    .D_N(_0836_),
    .X(_0847_));
 sky130_fd_sc_hd__o21a_4 _4289_ (.A1(_0704_),
    .A2(_0847_),
    .B1(_0803_),
    .X(_0858_));
 sky130_fd_sc_hd__o21ai_4 _4290_ (.A1(_0704_),
    .A2(_0847_),
    .B1(_0803_),
    .Y(_0869_));
 sky130_fd_sc_hd__nor2_2 _4291_ (.A(_0594_),
    .B(_0627_),
    .Y(_0880_));
 sky130_fd_sc_hd__o21ba_1 _4292_ (.A1(_0682_),
    .A2(_0880_),
    .B1_N(_0671_),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_4 _4293_ (.A0(_0726_),
    .A1(_0891_),
    .S(_0858_),
    .X(_0902_));
 sky130_fd_sc_hd__xnor2_4 _4294_ (.A(_0693_),
    .B(_0902_),
    .Y(_0913_));
 sky130_fd_sc_hd__xor2_4 _4295_ (.A(_0693_),
    .B(_0902_),
    .X(_0924_));
 sky130_fd_sc_hd__xnor2_4 _4296_ (.A(_0682_),
    .B(_0880_),
    .Y(_0935_));
 sky130_fd_sc_hd__o21a_2 _4297_ (.A1(_0616_),
    .A2(_0649_),
    .B1(_0869_),
    .X(_0946_));
 sky130_fd_sc_hd__xor2_4 _4298_ (.A(_0935_),
    .B(_0946_),
    .X(_0957_));
 sky130_fd_sc_hd__xnor2_4 _4299_ (.A(_0935_),
    .B(_0946_),
    .Y(_0968_));
 sky130_fd_sc_hd__and3_1 _4300_ (.A(net16),
    .B(_0154_),
    .C(_0616_),
    .X(_0979_));
 sky130_fd_sc_hd__or2_2 _4301_ (.A(_0627_),
    .B(_0979_),
    .X(_0990_));
 sky130_fd_sc_hd__nor2_1 _4302_ (.A(_0638_),
    .B(_0858_),
    .Y(_1001_));
 sky130_fd_sc_hd__xor2_4 _4303_ (.A(_0990_),
    .B(_1001_),
    .X(_1012_));
 sky130_fd_sc_hd__o2111ai_2 _4304_ (.A1(net19),
    .A2(_0165_),
    .B1(_0550_),
    .C1(_0561_),
    .D1(_0737_),
    .Y(_1023_));
 sky130_fd_sc_hd__a31o_1 _4305_ (.A1(_0517_),
    .A2(_0759_),
    .A3(_1023_),
    .B1(_0528_),
    .X(_1034_));
 sky130_fd_sc_hd__xnor2_1 _4306_ (.A(_0506_),
    .B(_1034_),
    .Y(_1045_));
 sky130_fd_sc_hd__xnor2_1 _4307_ (.A(_0792_),
    .B(_0836_),
    .Y(_1056_));
 sky130_fd_sc_hd__xnor2_1 _4308_ (.A(_0506_),
    .B(_0770_),
    .Y(_1067_));
 sky130_fd_sc_hd__a21o_1 _4309_ (.A1(_0869_),
    .A2(_1067_),
    .B1(_1056_),
    .X(_1078_));
 sky130_fd_sc_hd__nand2_1 _4310_ (.A(_1056_),
    .B(_1067_),
    .Y(_1089_));
 sky130_fd_sc_hd__o211a_4 _4311_ (.A1(_0858_),
    .A2(_1045_),
    .B1(_1078_),
    .C1(_1089_),
    .X(_1100_));
 sky130_fd_sc_hd__o22a_1 _4312_ (.A1(_0209_),
    .A2(_0297_),
    .B1(_0396_),
    .B2(_0429_),
    .X(_1111_));
 sky130_fd_sc_hd__and3_4 _4313_ (.A(_0176_),
    .B(_0209_),
    .C(_0429_),
    .X(_1122_));
 sky130_fd_sc_hd__and2_4 _4314_ (.A(_0814_),
    .B(_1122_),
    .X(_1133_));
 sky130_fd_sc_hd__nand2_8 _4315_ (.A(_0814_),
    .B(_1122_),
    .Y(_1144_));
 sky130_fd_sc_hd__or2_1 _4316_ (.A(net7),
    .B(_1133_),
    .X(_1155_));
 sky130_fd_sc_hd__o211a_1 _4317_ (.A1(net39),
    .A2(_1144_),
    .B1(_1155_),
    .C1(_1100_),
    .X(_1166_));
 sky130_fd_sc_hd__or2_1 _4318_ (.A(net6),
    .B(_1133_),
    .X(_1177_));
 sky130_fd_sc_hd__o211a_1 _4319_ (.A1(net38),
    .A2(_1144_),
    .B1(_1177_),
    .C1(_1100_),
    .X(_1188_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(_1166_),
    .A1(_1188_),
    .S(_0638_),
    .X(_1199_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(net5),
    .A1(net37),
    .S(_1133_),
    .X(_1210_));
 sky130_fd_sc_hd__mux2_1 _4322_ (.A0(net4),
    .A1(net36),
    .S(_1133_),
    .X(_1221_));
 sky130_fd_sc_hd__and2_1 _4323_ (.A(_1100_),
    .B(_1221_),
    .X(_1232_));
 sky130_fd_sc_hd__and3_1 _4324_ (.A(_0638_),
    .B(_1100_),
    .C(_1221_),
    .X(_1243_));
 sky130_fd_sc_hd__a31o_1 _4325_ (.A1(_0649_),
    .A2(_1100_),
    .A3(_1210_),
    .B1(_1243_),
    .X(_1254_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(_1199_),
    .A1(_1254_),
    .S(_1012_),
    .X(_1265_));
 sky130_fd_sc_hd__or2_1 _4327_ (.A(net31),
    .B(_1133_),
    .X(_1276_));
 sky130_fd_sc_hd__o211a_1 _4328_ (.A1(net63),
    .A2(_1144_),
    .B1(_1276_),
    .C1(_1100_),
    .X(_1287_));
 sky130_fd_sc_hd__or2_1 _4329_ (.A(net32),
    .B(_1133_),
    .X(_1298_));
 sky130_fd_sc_hd__o211a_1 _4330_ (.A1(net64),
    .A2(_1144_),
    .B1(_1298_),
    .C1(_1100_),
    .X(_1309_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(_1287_),
    .A1(_1309_),
    .S(_0649_),
    .X(_1320_));
 sky130_fd_sc_hd__nand2_1 _4332_ (.A(_0011_),
    .B(_1144_),
    .Y(_1331_));
 sky130_fd_sc_hd__o211a_1 _4333_ (.A1(net35),
    .A2(_1144_),
    .B1(_1331_),
    .C1(_1100_),
    .X(_1342_));
 sky130_fd_sc_hd__or2_1 _4334_ (.A(net2),
    .B(_1133_),
    .X(_1353_));
 sky130_fd_sc_hd__o211a_1 _4335_ (.A1(net34),
    .A2(_1144_),
    .B1(_1353_),
    .C1(_1100_),
    .X(_1364_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(_1342_),
    .A1(_1364_),
    .S(_0638_),
    .X(_1375_));
 sky130_fd_sc_hd__mux2_1 _4337_ (.A0(_1375_),
    .A1(_1320_),
    .S(_1012_),
    .X(_1386_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(_1265_),
    .A1(_1386_),
    .S(_0957_),
    .X(_1397_));
 sky130_fd_sc_hd__nand2_4 _4339_ (.A(_0704_),
    .B(_0814_),
    .Y(_1408_));
 sky130_fd_sc_hd__xnor2_4 _4340_ (.A(_0572_),
    .B(_0748_),
    .Y(_1419_));
 sky130_fd_sc_hd__xor2_4 _4341_ (.A(_1408_),
    .B(_1419_),
    .X(_1430_));
 sky130_fd_sc_hd__xnor2_4 _4342_ (.A(_1408_),
    .B(_1419_),
    .Y(_1441_));
 sky130_fd_sc_hd__mux2_1 _4343_ (.A0(net29),
    .A1(net61),
    .S(_1133_),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _4344_ (.A0(net30),
    .A1(net62),
    .S(_1133_),
    .X(_1463_));
 sky130_fd_sc_hd__and2_1 _4345_ (.A(_1100_),
    .B(_1463_),
    .X(_1474_));
 sky130_fd_sc_hd__and3_1 _4346_ (.A(_0649_),
    .B(_1100_),
    .C(_1463_),
    .X(_1485_));
 sky130_fd_sc_hd__a31o_1 _4347_ (.A1(_0638_),
    .A2(_1100_),
    .A3(_1452_),
    .B1(_1485_),
    .X(_1496_));
 sky130_fd_sc_hd__mux2_1 _4348_ (.A0(net27),
    .A1(net59),
    .S(_1133_),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _4349_ (.A0(net28),
    .A1(net60),
    .S(_1133_),
    .X(_1518_));
 sky130_fd_sc_hd__or2_1 _4350_ (.A(_0638_),
    .B(_1518_),
    .X(_1529_));
 sky130_fd_sc_hd__o211a_1 _4351_ (.A1(_0649_),
    .A2(_1507_),
    .B1(_1529_),
    .C1(_1100_),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_1 _4352_ (.A0(_1496_),
    .A1(_1540_),
    .S(_1012_),
    .X(_1551_));
 sky130_fd_sc_hd__mux4_1 _4353_ (.A0(net26),
    .A1(net23),
    .A2(net58),
    .A3(net55),
    .S0(_0638_),
    .S1(_1133_),
    .X(_1562_));
 sky130_fd_sc_hd__nand2_1 _4354_ (.A(_1100_),
    .B(_1562_),
    .Y(_1573_));
 sky130_fd_sc_hd__nor2_1 _4355_ (.A(_1012_),
    .B(_1573_),
    .Y(_1584_));
 sky130_fd_sc_hd__mux4_1 _4356_ (.A0(net44),
    .A1(net33),
    .A2(net12),
    .A3(net1),
    .S0(_0638_),
    .S1(_1144_),
    .X(_1595_));
 sky130_fd_sc_hd__a31o_1 _4357_ (.A1(_1012_),
    .A2(_1100_),
    .A3(_1595_),
    .B1(_0968_),
    .X(_1606_));
 sky130_fd_sc_hd__o221a_1 _4358_ (.A1(_0957_),
    .A2(_1551_),
    .B1(_1584_),
    .B2(_1606_),
    .C1(_0913_),
    .X(_1617_));
 sky130_fd_sc_hd__a211o_1 _4359_ (.A1(_0924_),
    .A2(_1397_),
    .B1(_1430_),
    .C1(_1617_),
    .X(_1628_));
 sky130_fd_sc_hd__nor2_1 _4360_ (.A(_0759_),
    .B(_0869_),
    .Y(_1639_));
 sky130_fd_sc_hd__a31o_1 _4361_ (.A1(_0561_),
    .A2(_0869_),
    .A3(_1023_),
    .B1(_1639_),
    .X(_1650_));
 sky130_fd_sc_hd__xor2_4 _4362_ (.A(_0825_),
    .B(_1650_),
    .X(_1661_));
 sky130_fd_sc_hd__nor2_4 _4363_ (.A(_1430_),
    .B(_1661_),
    .Y(_1672_));
 sky130_fd_sc_hd__or2_1 _4364_ (.A(_1430_),
    .B(_1661_),
    .X(_1683_));
 sky130_fd_sc_hd__or4_1 _4365_ (.A(net19),
    .B(net21),
    .C(net22),
    .D(net24),
    .X(_1694_));
 sky130_fd_sc_hd__or4_1 _4366_ (.A(net16),
    .B(net18),
    .C(net17),
    .D(net20),
    .X(_1705_));
 sky130_fd_sc_hd__or2_4 _4367_ (.A(_1694_),
    .B(_1705_),
    .X(_1716_));
 sky130_fd_sc_hd__inv_2 _4368_ (.A(_1716_),
    .Y(_1727_));
 sky130_fd_sc_hd__or4_1 _4369_ (.A(net51),
    .B(net54),
    .C(net53),
    .D(net56),
    .X(_1738_));
 sky130_fd_sc_hd__or4_1 _4370_ (.A(net48),
    .B(net50),
    .C(net49),
    .D(net52),
    .X(_1749_));
 sky130_fd_sc_hd__or2_4 _4371_ (.A(_1738_),
    .B(_1749_),
    .X(_1760_));
 sky130_fd_sc_hd__inv_2 _4372_ (.A(_1760_),
    .Y(_1771_));
 sky130_fd_sc_hd__o211a_1 _4373_ (.A1(_1144_),
    .A2(_1760_),
    .B1(_1716_),
    .C1(_1100_),
    .X(_1782_));
 sky130_fd_sc_hd__or2_1 _4374_ (.A(net15),
    .B(_1133_),
    .X(_1793_));
 sky130_fd_sc_hd__o211a_1 _4375_ (.A1(net47),
    .A2(_1144_),
    .B1(_1793_),
    .C1(_1100_),
    .X(_1804_));
 sky130_fd_sc_hd__mux2_1 _4376_ (.A0(_1782_),
    .A1(_1804_),
    .S(_0638_),
    .X(_1815_));
 sky130_fd_sc_hd__or2_1 _4377_ (.A(net14),
    .B(_1133_),
    .X(_1826_));
 sky130_fd_sc_hd__o211a_1 _4378_ (.A1(net46),
    .A2(_1144_),
    .B1(_1826_),
    .C1(_1100_),
    .X(_1837_));
 sky130_fd_sc_hd__nand2_1 _4379_ (.A(_0000_),
    .B(_1144_),
    .Y(_1848_));
 sky130_fd_sc_hd__o211a_1 _4380_ (.A1(net45),
    .A2(_1144_),
    .B1(_1848_),
    .C1(_1100_),
    .X(_1859_));
 sky130_fd_sc_hd__mux2_1 _4381_ (.A0(_1837_),
    .A1(_1859_),
    .S(_0638_),
    .X(_1870_));
 sky130_fd_sc_hd__mux2_1 _4382_ (.A0(_1815_),
    .A1(_1870_),
    .S(_1012_),
    .X(_1881_));
 sky130_fd_sc_hd__or2_1 _4383_ (.A(net11),
    .B(_1133_),
    .X(_1892_));
 sky130_fd_sc_hd__o211a_1 _4384_ (.A1(net43),
    .A2(_1144_),
    .B1(_1892_),
    .C1(_1100_),
    .X(_1903_));
 sky130_fd_sc_hd__or2_1 _4385_ (.A(net10),
    .B(_1133_),
    .X(_1914_));
 sky130_fd_sc_hd__o211a_1 _4386_ (.A1(net42),
    .A2(_1144_),
    .B1(_1914_),
    .C1(_1100_),
    .X(_1925_));
 sky130_fd_sc_hd__mux2_1 _4387_ (.A0(_1903_),
    .A1(_1925_),
    .S(_0638_),
    .X(_1936_));
 sky130_fd_sc_hd__or2_1 _4388_ (.A(net9),
    .B(_1133_),
    .X(_1947_));
 sky130_fd_sc_hd__o211a_1 _4389_ (.A1(net41),
    .A2(_1144_),
    .B1(_1947_),
    .C1(_1100_),
    .X(_1958_));
 sky130_fd_sc_hd__or2_1 _4390_ (.A(net8),
    .B(_1133_),
    .X(_1969_));
 sky130_fd_sc_hd__o211a_1 _4391_ (.A1(net40),
    .A2(_1144_),
    .B1(_1969_),
    .C1(_1100_),
    .X(_1980_));
 sky130_fd_sc_hd__mux2_1 _4392_ (.A0(_1958_),
    .A1(_1980_),
    .S(_0638_),
    .X(_1991_));
 sky130_fd_sc_hd__mux2_1 _4393_ (.A0(_1936_),
    .A1(_1991_),
    .S(_1012_),
    .X(_2002_));
 sky130_fd_sc_hd__mux2_1 _4394_ (.A0(_1881_),
    .A1(_2002_),
    .S(_0957_),
    .X(_2013_));
 sky130_fd_sc_hd__nor2_1 _4395_ (.A(_0924_),
    .B(_1661_),
    .Y(_2024_));
 sky130_fd_sc_hd__or2_1 _4396_ (.A(_0924_),
    .B(_1661_),
    .X(_2035_));
 sky130_fd_sc_hd__a21o_1 _4397_ (.A1(_2013_),
    .A2(_2024_),
    .B1(_1672_),
    .X(_2046_));
 sky130_fd_sc_hd__and2_1 _4398_ (.A(_1628_),
    .B(_2046_),
    .X(_2057_));
 sky130_fd_sc_hd__mux2_1 _4399_ (.A0(net33),
    .A1(_2057_),
    .S(_0814_),
    .X(_2068_));
 sky130_fd_sc_hd__mux2_1 _4400_ (.A0(net1),
    .A1(_2057_),
    .S(_0858_),
    .X(_2079_));
 sky130_fd_sc_hd__nand2_1 _4401_ (.A(_2068_),
    .B(_2079_),
    .Y(_2090_));
 sky130_fd_sc_hd__and2_1 _4402_ (.A(_0638_),
    .B(_1782_),
    .X(_2101_));
 sky130_fd_sc_hd__nand2_1 _4403_ (.A(_0990_),
    .B(_2101_),
    .Y(_2112_));
 sky130_fd_sc_hd__inv_2 _4404_ (.A(_2112_),
    .Y(_2123_));
 sky130_fd_sc_hd__mux2_1 _4405_ (.A0(_1804_),
    .A1(_1837_),
    .S(_0638_),
    .X(_2134_));
 sky130_fd_sc_hd__mux2_1 _4406_ (.A0(_1859_),
    .A1(_1903_),
    .S(_0638_),
    .X(_2145_));
 sky130_fd_sc_hd__mux2_1 _4407_ (.A0(_2134_),
    .A1(_2145_),
    .S(_1012_),
    .X(_2156_));
 sky130_fd_sc_hd__mux2_1 _4408_ (.A0(_2123_),
    .A1(_2156_),
    .S(_0957_),
    .X(_2167_));
 sky130_fd_sc_hd__and3_1 _4409_ (.A(_0913_),
    .B(_1672_),
    .C(_2167_),
    .X(_2178_));
 sky130_fd_sc_hd__mux2_1 _4410_ (.A0(net43),
    .A1(_2178_),
    .S(net98),
    .X(_2189_));
 sky130_fd_sc_hd__mux2_1 _4411_ (.A0(net11),
    .A1(_2178_),
    .S(_0858_),
    .X(_2200_));
 sky130_fd_sc_hd__nand2b_1 _4412_ (.A_N(_2189_),
    .B(_2200_),
    .Y(_2211_));
 sky130_fd_sc_hd__nand2_1 _4413_ (.A(_1012_),
    .B(_1815_),
    .Y(_2222_));
 sky130_fd_sc_hd__mux2_1 _4414_ (.A0(_1870_),
    .A1(_1936_),
    .S(_1012_),
    .X(_2233_));
 sky130_fd_sc_hd__inv_2 _4415_ (.A(_2233_),
    .Y(_2244_));
 sky130_fd_sc_hd__mux2_1 _4416_ (.A0(_2222_),
    .A1(_2244_),
    .S(_0957_),
    .X(_2255_));
 sky130_fd_sc_hd__nor2_1 _4417_ (.A(_2035_),
    .B(_2255_),
    .Y(_2266_));
 sky130_fd_sc_hd__and2_1 _4418_ (.A(_1441_),
    .B(_2266_),
    .X(_2277_));
 sky130_fd_sc_hd__mux2_1 _4419_ (.A0(net42),
    .A1(_2277_),
    .S(net98),
    .X(_2288_));
 sky130_fd_sc_hd__mux2_1 _4420_ (.A0(net10),
    .A1(_2277_),
    .S(_0858_),
    .X(_2299_));
 sky130_fd_sc_hd__mux2_1 _4421_ (.A0(_2101_),
    .A1(_2134_),
    .S(_1012_),
    .X(_2310_));
 sky130_fd_sc_hd__mux2_1 _4422_ (.A0(_1925_),
    .A1(_1958_),
    .S(_0638_),
    .X(_2321_));
 sky130_fd_sc_hd__mux2_1 _4423_ (.A0(_2145_),
    .A1(_2321_),
    .S(_1012_),
    .X(_2332_));
 sky130_fd_sc_hd__inv_2 _4424_ (.A(_2332_),
    .Y(_2343_));
 sky130_fd_sc_hd__mux2_1 _4425_ (.A0(_2310_),
    .A1(_2332_),
    .S(_0957_),
    .X(_2354_));
 sky130_fd_sc_hd__and3_1 _4426_ (.A(_0913_),
    .B(_1672_),
    .C(_2354_),
    .X(_2365_));
 sky130_fd_sc_hd__mux2_1 _4427_ (.A0(net41),
    .A1(_2365_),
    .S(net98),
    .X(_2376_));
 sky130_fd_sc_hd__mux2_1 _4428_ (.A0(net9),
    .A1(_2365_),
    .S(_0858_),
    .X(_2387_));
 sky130_fd_sc_hd__inv_2 _4429_ (.A(_2387_),
    .Y(_2398_));
 sky130_fd_sc_hd__xnor2_1 _4430_ (.A(_2288_),
    .B(_2299_),
    .Y(_2409_));
 sky130_fd_sc_hd__o211a_1 _4431_ (.A1(_2376_),
    .A2(_2398_),
    .B1(_2409_),
    .C1(_2211_),
    .X(_2420_));
 sky130_fd_sc_hd__nand2_1 _4432_ (.A(_0957_),
    .B(_2310_),
    .Y(_2431_));
 sky130_fd_sc_hd__nor2_1 _4433_ (.A(_2035_),
    .B(_2431_),
    .Y(_2442_));
 sky130_fd_sc_hd__and2_1 _4434_ (.A(_1441_),
    .B(_2442_),
    .X(_2453_));
 sky130_fd_sc_hd__mux2_1 _4435_ (.A0(net46),
    .A1(_2453_),
    .S(net98),
    .X(_2464_));
 sky130_fd_sc_hd__mux2_1 _4436_ (.A0(net14),
    .A1(_2453_),
    .S(_0858_),
    .X(_2475_));
 sky130_fd_sc_hd__inv_2 _4437_ (.A(_2475_),
    .Y(_2486_));
 sky130_fd_sc_hd__nand2_1 _4438_ (.A(_0957_),
    .B(_1881_),
    .Y(_2497_));
 sky130_fd_sc_hd__or2_1 _4439_ (.A(_2035_),
    .B(_2497_),
    .X(_2508_));
 sky130_fd_sc_hd__nor2_1 _4440_ (.A(_1430_),
    .B(_2508_),
    .Y(_2519_));
 sky130_fd_sc_hd__mux2_1 _4441_ (.A0(net45),
    .A1(_2519_),
    .S(net98),
    .X(_2530_));
 sky130_fd_sc_hd__mux2_1 _4442_ (.A0(net13),
    .A1(_2519_),
    .S(_0858_),
    .X(_2541_));
 sky130_fd_sc_hd__inv_2 _4443_ (.A(_2541_),
    .Y(_2552_));
 sky130_fd_sc_hd__a22o_1 _4444_ (.A1(_2464_),
    .A2(_2486_),
    .B1(_2530_),
    .B2(_2552_),
    .X(_2563_));
 sky130_fd_sc_hd__and2b_1 _4445_ (.A_N(_2200_),
    .B(_2189_),
    .X(_2574_));
 sky130_fd_sc_hd__nor2_1 _4446_ (.A(_0968_),
    .B(_2222_),
    .Y(_2585_));
 sky130_fd_sc_hd__nand2_1 _4447_ (.A(_2024_),
    .B(_2585_),
    .Y(_2596_));
 sky130_fd_sc_hd__nor2_1 _4448_ (.A(_1430_),
    .B(_2596_),
    .Y(_2607_));
 sky130_fd_sc_hd__mux2_1 _4449_ (.A0(net15),
    .A1(_2607_),
    .S(_0858_),
    .X(_2618_));
 sky130_fd_sc_hd__inv_2 _4450_ (.A(_2618_),
    .Y(_2629_));
 sky130_fd_sc_hd__o22a_1 _4451_ (.A1(_2464_),
    .A2(_2486_),
    .B1(_2629_),
    .B2(net47),
    .X(_2640_));
 sky130_fd_sc_hd__and3_1 _4452_ (.A(_0913_),
    .B(_1672_),
    .C(_2013_),
    .X(_2651_));
 sky130_fd_sc_hd__mux2_1 _4453_ (.A0(net40),
    .A1(_2651_),
    .S(net98),
    .X(_2662_));
 sky130_fd_sc_hd__mux2_1 _4454_ (.A0(net8),
    .A1(_2651_),
    .S(_0858_),
    .X(_2673_));
 sky130_fd_sc_hd__inv_2 _4455_ (.A(_2673_),
    .Y(_2684_));
 sky130_fd_sc_hd__a22o_1 _4456_ (.A1(_2376_),
    .A2(_2398_),
    .B1(_2662_),
    .B2(_2684_),
    .X(_2695_));
 sky130_fd_sc_hd__or2_1 _4457_ (.A(_2530_),
    .B(_2552_),
    .X(_2706_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(net47),
    .A1(_2607_),
    .S(net98),
    .X(_2717_));
 sky130_fd_sc_hd__a21o_1 _4459_ (.A1(_2629_),
    .A2(_2717_),
    .B1(_0858_),
    .X(_2728_));
 sky130_fd_sc_hd__and3b_1 _4460_ (.A_N(_2728_),
    .B(_2640_),
    .C(_0803_),
    .X(_2739_));
 sky130_fd_sc_hd__o21ai_1 _4461_ (.A1(_2662_),
    .A2(_2684_),
    .B1(_2706_),
    .Y(_2750_));
 sky130_fd_sc_hd__nand2_1 _4462_ (.A(_2420_),
    .B(_2739_),
    .Y(_2761_));
 sky130_fd_sc_hd__or4_1 _4463_ (.A(_2563_),
    .B(_2574_),
    .C(_2750_),
    .D(_2761_),
    .X(_2772_));
 sky130_fd_sc_hd__nor2_1 _4464_ (.A(_2695_),
    .B(_2772_),
    .Y(_2783_));
 sky130_fd_sc_hd__inv_2 _4465_ (.A(_2783_),
    .Y(_2794_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(_1166_),
    .A1(_1980_),
    .S(_0649_),
    .X(_2805_));
 sky130_fd_sc_hd__mux2_1 _4467_ (.A0(_2321_),
    .A1(_2805_),
    .S(_1012_),
    .X(_2816_));
 sky130_fd_sc_hd__inv_2 _4468_ (.A(_2816_),
    .Y(_2827_));
 sky130_fd_sc_hd__mux2_1 _4469_ (.A0(_2156_),
    .A1(_2816_),
    .S(_0957_),
    .X(_2838_));
 sky130_fd_sc_hd__or2_1 _4470_ (.A(_0924_),
    .B(_2838_),
    .X(_2849_));
 sky130_fd_sc_hd__nor2_1 _4471_ (.A(_0968_),
    .B(_2112_),
    .Y(_2860_));
 sky130_fd_sc_hd__o211a_1 _4472_ (.A1(_0913_),
    .A2(_2860_),
    .B1(_2849_),
    .C1(_1672_),
    .X(_2871_));
 sky130_fd_sc_hd__inv_2 _4473_ (.A(_2871_),
    .Y(_2882_));
 sky130_fd_sc_hd__mux2_1 _4474_ (.A0(_0088_),
    .A1(_2882_),
    .S(net98),
    .X(_2893_));
 sky130_fd_sc_hd__mux2_1 _4475_ (.A0(net39),
    .A1(_2871_),
    .S(net98),
    .X(_2904_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(net7),
    .A1(_2871_),
    .S(_0858_),
    .X(_2915_));
 sky130_fd_sc_hd__nand2_1 _4477_ (.A(_2893_),
    .B(_2915_),
    .Y(_2926_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(_1991_),
    .A1(_1199_),
    .S(_1012_),
    .X(_2937_));
 sky130_fd_sc_hd__inv_2 _4479_ (.A(_2937_),
    .Y(_2948_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(_2244_),
    .A1(_2948_),
    .S(_0957_),
    .X(_2959_));
 sky130_fd_sc_hd__nand2_1 _4481_ (.A(_0913_),
    .B(_2959_),
    .Y(_2970_));
 sky130_fd_sc_hd__o211a_1 _4482_ (.A1(_0913_),
    .A2(_2585_),
    .B1(_2970_),
    .C1(_1672_),
    .X(_2981_));
 sky130_fd_sc_hd__mux2_1 _4483_ (.A0(net38),
    .A1(_2981_),
    .S(net98),
    .X(_2992_));
 sky130_fd_sc_hd__mux2_1 _4484_ (.A0(net6),
    .A1(_2981_),
    .S(_0858_),
    .X(_3003_));
 sky130_fd_sc_hd__inv_2 _4485_ (.A(_3003_),
    .Y(_3014_));
 sky130_fd_sc_hd__a2bb2o_1 _4486_ (.A1_N(_2893_),
    .A2_N(_2915_),
    .B1(_2992_),
    .B2(_3014_),
    .X(_3025_));
 sky130_fd_sc_hd__and3_1 _4487_ (.A(_0638_),
    .B(_1100_),
    .C(_1210_),
    .X(_3036_));
 sky130_fd_sc_hd__a21oi_1 _4488_ (.A1(_0649_),
    .A2(_1188_),
    .B1(_3036_),
    .Y(_3047_));
 sky130_fd_sc_hd__mux2_1 _4489_ (.A0(_1232_),
    .A1(_1342_),
    .S(_0638_),
    .X(_3058_));
 sky130_fd_sc_hd__inv_2 _4490_ (.A(_3058_),
    .Y(_3069_));
 sky130_fd_sc_hd__mux2_1 _4491_ (.A0(_3047_),
    .A1(_3069_),
    .S(_1012_),
    .X(_3080_));
 sky130_fd_sc_hd__mux2_1 _4492_ (.A0(_2827_),
    .A1(_3080_),
    .S(_0957_),
    .X(_3091_));
 sky130_fd_sc_hd__nand2_1 _4493_ (.A(_0913_),
    .B(_3091_),
    .Y(_3102_));
 sky130_fd_sc_hd__o211a_1 _4494_ (.A1(_0913_),
    .A2(_2167_),
    .B1(_3102_),
    .C1(_1672_),
    .X(_3113_));
 sky130_fd_sc_hd__mux2_1 _4495_ (.A0(net35),
    .A1(_3113_),
    .S(net98),
    .X(_3124_));
 sky130_fd_sc_hd__inv_2 _4496_ (.A(_3124_),
    .Y(_3135_));
 sky130_fd_sc_hd__mux2_1 _4497_ (.A0(net3),
    .A1(_3113_),
    .S(_0858_),
    .X(_3146_));
 sky130_fd_sc_hd__mux2_1 _4498_ (.A0(_1265_),
    .A1(_2002_),
    .S(_0968_),
    .X(_3157_));
 sky130_fd_sc_hd__nand2_1 _4499_ (.A(_0924_),
    .B(_2497_),
    .Y(_3168_));
 sky130_fd_sc_hd__o211a_1 _4500_ (.A1(_0924_),
    .A2(_3157_),
    .B1(_3168_),
    .C1(_1672_),
    .X(_3179_));
 sky130_fd_sc_hd__inv_2 _4501_ (.A(_3179_),
    .Y(_3190_));
 sky130_fd_sc_hd__mux2_1 _4502_ (.A0(_0066_),
    .A1(_3190_),
    .S(net98),
    .X(_3201_));
 sky130_fd_sc_hd__mux2_1 _4503_ (.A0(net36),
    .A1(_3179_),
    .S(net98),
    .X(_3212_));
 sky130_fd_sc_hd__mux2_1 _4504_ (.A0(net4),
    .A1(_3179_),
    .S(_0858_),
    .X(_3223_));
 sky130_fd_sc_hd__nor2_1 _4505_ (.A(_1012_),
    .B(_2805_),
    .Y(_3234_));
 sky130_fd_sc_hd__a21o_1 _4506_ (.A1(_1012_),
    .A2(_3047_),
    .B1(_3234_),
    .X(_3245_));
 sky130_fd_sc_hd__mux2_1 _4507_ (.A0(_2343_),
    .A1(_3245_),
    .S(_0957_),
    .X(_3256_));
 sky130_fd_sc_hd__a21o_1 _4508_ (.A1(_0924_),
    .A2(_2431_),
    .B1(_1683_),
    .X(_3267_));
 sky130_fd_sc_hd__a21oi_2 _4509_ (.A1(_0913_),
    .A2(_3256_),
    .B1(_3267_),
    .Y(_3278_));
 sky130_fd_sc_hd__inv_2 _4510_ (.A(_3278_),
    .Y(_3289_));
 sky130_fd_sc_hd__mux2_1 _4511_ (.A0(_0077_),
    .A1(_3289_),
    .S(net98),
    .X(_3300_));
 sky130_fd_sc_hd__mux2_1 _4512_ (.A0(net37),
    .A1(_3278_),
    .S(net98),
    .X(_3311_));
 sky130_fd_sc_hd__mux2_1 _4513_ (.A0(net5),
    .A1(_3278_),
    .S(_0858_),
    .X(_3322_));
 sky130_fd_sc_hd__a22o_1 _4514_ (.A1(_3201_),
    .A2(_3223_),
    .B1(_3300_),
    .B2(_3322_),
    .X(_3333_));
 sky130_fd_sc_hd__mux2_1 _4515_ (.A0(_1254_),
    .A1(_1375_),
    .S(_1012_),
    .X(_3344_));
 sky130_fd_sc_hd__mux2_1 _4516_ (.A0(_2937_),
    .A1(_3344_),
    .S(_0957_),
    .X(_3355_));
 sky130_fd_sc_hd__nand2_1 _4517_ (.A(_0924_),
    .B(_2255_),
    .Y(_3365_));
 sky130_fd_sc_hd__o211a_1 _4518_ (.A1(_0924_),
    .A2(_3355_),
    .B1(_3365_),
    .C1(_1672_),
    .X(_3375_));
 sky130_fd_sc_hd__mux2_1 _4519_ (.A0(net34),
    .A1(_3375_),
    .S(net98),
    .X(_3386_));
 sky130_fd_sc_hd__inv_2 _4520_ (.A(_3386_),
    .Y(_3397_));
 sky130_fd_sc_hd__mux2_1 _4521_ (.A0(net2),
    .A1(_3375_),
    .S(_0858_),
    .X(_3408_));
 sky130_fd_sc_hd__a221o_1 _4522_ (.A1(_3135_),
    .A2(_3146_),
    .B1(_3397_),
    .B2(_3408_),
    .C1(_3333_),
    .X(_3419_));
 sky130_fd_sc_hd__mux2_1 _4523_ (.A0(_1309_),
    .A1(_1364_),
    .S(_0649_),
    .X(_3429_));
 sky130_fd_sc_hd__mux2_1 _4524_ (.A0(_3058_),
    .A1(_3429_),
    .S(_1012_),
    .X(_3438_));
 sky130_fd_sc_hd__nand2_1 _4525_ (.A(_0957_),
    .B(_3438_),
    .Y(_3448_));
 sky130_fd_sc_hd__o21ai_1 _4526_ (.A1(_0957_),
    .A2(_3245_),
    .B1(_3448_),
    .Y(_3457_));
 sky130_fd_sc_hd__or2_1 _4527_ (.A(_0913_),
    .B(_2354_),
    .X(_3467_));
 sky130_fd_sc_hd__o211a_1 _4528_ (.A1(_0924_),
    .A2(_3457_),
    .B1(_3467_),
    .C1(_1672_),
    .X(_3477_));
 sky130_fd_sc_hd__inv_2 _4529_ (.A(_3477_),
    .Y(_3486_));
 sky130_fd_sc_hd__mux2_1 _4530_ (.A0(_0044_),
    .A1(_3486_),
    .S(net98),
    .X(_3496_));
 sky130_fd_sc_hd__mux2_1 _4531_ (.A0(net64),
    .A1(_3477_),
    .S(net98),
    .X(_3505_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(net32),
    .A1(_3477_),
    .S(_0858_),
    .X(_3515_));
 sky130_fd_sc_hd__o22a_1 _4533_ (.A1(_3397_),
    .A2(_3408_),
    .B1(_3496_),
    .B2(_3515_),
    .X(_3524_));
 sky130_fd_sc_hd__and2_1 _4534_ (.A(_3496_),
    .B(_3515_),
    .X(_3534_));
 sky130_fd_sc_hd__or2_1 _4535_ (.A(_0924_),
    .B(_1397_),
    .X(_3544_));
 sky130_fd_sc_hd__o211a_1 _4536_ (.A1(_0913_),
    .A2(_2013_),
    .B1(_3544_),
    .C1(_1672_),
    .X(_3553_));
 sky130_fd_sc_hd__mux2_1 _4537_ (.A0(net63),
    .A1(_3553_),
    .S(net98),
    .X(_3563_));
 sky130_fd_sc_hd__mux2_1 _4538_ (.A0(net31),
    .A1(_3553_),
    .S(_0858_),
    .X(_3573_));
 sky130_fd_sc_hd__or3b_1 _4539_ (.A(_3534_),
    .B(_3573_),
    .C_N(_3563_),
    .X(_3583_));
 sky130_fd_sc_hd__a21o_1 _4540_ (.A1(_3524_),
    .A2(_3583_),
    .B1(_3419_),
    .X(_3593_));
 sky130_fd_sc_hd__or2_1 _4541_ (.A(_3300_),
    .B(_3322_),
    .X(_3603_));
 sky130_fd_sc_hd__o22a_1 _4542_ (.A1(_3135_),
    .A2(_3146_),
    .B1(_3201_),
    .B2(_3223_),
    .X(_3613_));
 sky130_fd_sc_hd__o21a_1 _4543_ (.A1(_3333_),
    .A2(_3613_),
    .B1(_3603_),
    .X(_3623_));
 sky130_fd_sc_hd__a2bb2o_1 _4544_ (.A1_N(_2992_),
    .A2_N(_3014_),
    .B1(_3593_),
    .B2(_3623_),
    .X(_3633_));
 sky130_fd_sc_hd__nand2b_1 _4545_ (.A_N(_3025_),
    .B(_3633_),
    .Y(_3641_));
 sky130_fd_sc_hd__nor2_1 _4546_ (.A(_0957_),
    .B(_3344_),
    .Y(_3642_));
 sky130_fd_sc_hd__mux2_1 _4547_ (.A0(_1320_),
    .A1(_1496_),
    .S(_1012_),
    .X(_3643_));
 sky130_fd_sc_hd__o21ai_1 _4548_ (.A1(_0968_),
    .A2(_3643_),
    .B1(_0913_),
    .Y(_3644_));
 sky130_fd_sc_hd__o221a_1 _4549_ (.A1(_0913_),
    .A2(_2959_),
    .B1(_3642_),
    .B2(_3644_),
    .C1(_1441_),
    .X(_3645_));
 sky130_fd_sc_hd__a21oi_1 _4550_ (.A1(_1683_),
    .A2(_2596_),
    .B1(_3645_),
    .Y(_3646_));
 sky130_fd_sc_hd__mux2_1 _4551_ (.A0(net61),
    .A1(_3646_),
    .S(net98),
    .X(_3647_));
 sky130_fd_sc_hd__mux2_1 _4552_ (.A0(net29),
    .A1(_3646_),
    .S(_0858_),
    .X(_3648_));
 sky130_fd_sc_hd__inv_2 _4553_ (.A(_3648_),
    .Y(_3649_));
 sky130_fd_sc_hd__nand2_1 _4554_ (.A(_0924_),
    .B(_2838_),
    .Y(_3650_));
 sky130_fd_sc_hd__and2b_1 _4555_ (.A_N(_1012_),
    .B(_3429_),
    .X(_3651_));
 sky130_fd_sc_hd__mux2_1 _4556_ (.A0(_1287_),
    .A1(_1474_),
    .S(_0638_),
    .X(_3652_));
 sky130_fd_sc_hd__a21oi_1 _4557_ (.A1(_1012_),
    .A2(_3652_),
    .B1(_3651_),
    .Y(_3653_));
 sky130_fd_sc_hd__mux2_1 _4558_ (.A0(_3080_),
    .A1(_3653_),
    .S(_0957_),
    .X(_3654_));
 sky130_fd_sc_hd__o211a_1 _4559_ (.A1(_0924_),
    .A2(_3654_),
    .B1(_3650_),
    .C1(_1441_),
    .X(_3655_));
 sky130_fd_sc_hd__nand2_1 _4560_ (.A(_2024_),
    .B(_2860_),
    .Y(_3656_));
 sky130_fd_sc_hd__a21oi_1 _4561_ (.A1(_1683_),
    .A2(_3656_),
    .B1(_3655_),
    .Y(_3657_));
 sky130_fd_sc_hd__mux2_1 _4562_ (.A0(net62),
    .A1(_3657_),
    .S(net98),
    .X(_3658_));
 sky130_fd_sc_hd__and2_1 _4563_ (.A(_0858_),
    .B(_3657_),
    .X(_3659_));
 sky130_fd_sc_hd__a21oi_1 _4564_ (.A1(net30),
    .A2(_0869_),
    .B1(_3659_),
    .Y(_3660_));
 sky130_fd_sc_hd__a21o_1 _4565_ (.A1(net30),
    .A2(_0869_),
    .B1(_3659_),
    .X(_3661_));
 sky130_fd_sc_hd__a22o_1 _4566_ (.A1(_3647_),
    .A2(_3649_),
    .B1(_3658_),
    .B2(_3660_),
    .X(_3662_));
 sky130_fd_sc_hd__inv_2 _4567_ (.A(_3662_),
    .Y(_3663_));
 sky130_fd_sc_hd__nand2_1 _4568_ (.A(_0924_),
    .B(_3157_),
    .Y(_3664_));
 sky130_fd_sc_hd__o21a_1 _4569_ (.A1(_0957_),
    .A2(_1386_),
    .B1(_0913_),
    .X(_3665_));
 sky130_fd_sc_hd__o21ai_1 _4570_ (.A1(_0968_),
    .A2(_1551_),
    .B1(_3665_),
    .Y(_3666_));
 sky130_fd_sc_hd__a32o_1 _4571_ (.A1(_1441_),
    .A2(_3664_),
    .A3(_3666_),
    .B1(_1683_),
    .B2(_2508_),
    .X(_3667_));
 sky130_fd_sc_hd__inv_2 _4572_ (.A(_3667_),
    .Y(_3668_));
 sky130_fd_sc_hd__mux2_1 _4573_ (.A0(net59),
    .A1(_3668_),
    .S(net98),
    .X(_3669_));
 sky130_fd_sc_hd__mux2_1 _4574_ (.A0(_4187_),
    .A1(_3667_),
    .S(_0858_),
    .X(_3670_));
 sky130_fd_sc_hd__inv_2 _4575_ (.A(_3670_),
    .Y(_3671_));
 sky130_fd_sc_hd__nor2_1 _4576_ (.A(_0033_),
    .B(net98),
    .Y(_3672_));
 sky130_fd_sc_hd__or2_1 _4577_ (.A(_0638_),
    .B(_1452_),
    .X(_3673_));
 sky130_fd_sc_hd__o211a_1 _4578_ (.A1(_0649_),
    .A2(_1518_),
    .B1(_3673_),
    .C1(_1100_),
    .X(_3674_));
 sky130_fd_sc_hd__inv_2 _4579_ (.A(_3674_),
    .Y(_3675_));
 sky130_fd_sc_hd__mux2_1 _4580_ (.A0(_3652_),
    .A1(_3674_),
    .S(_1012_),
    .X(_3676_));
 sky130_fd_sc_hd__mux2_1 _4581_ (.A0(_3438_),
    .A1(_3676_),
    .S(_0957_),
    .X(_3677_));
 sky130_fd_sc_hd__nand2_1 _4582_ (.A(_0913_),
    .B(_3677_),
    .Y(_3678_));
 sky130_fd_sc_hd__o21ai_1 _4583_ (.A1(_0913_),
    .A2(_3256_),
    .B1(_3678_),
    .Y(_3679_));
 sky130_fd_sc_hd__o22a_1 _4584_ (.A1(_1672_),
    .A2(_2442_),
    .B1(_3679_),
    .B2(_1430_),
    .X(_3680_));
 sky130_fd_sc_hd__a21oi_1 _4585_ (.A1(net98),
    .A2(_3680_),
    .B1(_3672_),
    .Y(_3681_));
 sky130_fd_sc_hd__inv_2 _4586_ (.A(_3681_),
    .Y(_3682_));
 sky130_fd_sc_hd__mux2_1 _4587_ (.A0(net28),
    .A1(_3680_),
    .S(_0858_),
    .X(_3683_));
 sky130_fd_sc_hd__inv_2 _4588_ (.A(_3683_),
    .Y(_3684_));
 sky130_fd_sc_hd__a221o_1 _4589_ (.A1(_3669_),
    .A2(_3670_),
    .B1(_3682_),
    .B2(_3684_),
    .C1(_3662_),
    .X(_3685_));
 sky130_fd_sc_hd__nor2_1 _4590_ (.A(_3669_),
    .B(_3670_),
    .Y(_3686_));
 sky130_fd_sc_hd__mux4_1 _4591_ (.A0(net27),
    .A1(net26),
    .A2(net59),
    .A3(net58),
    .S0(_0638_),
    .S1(_1133_),
    .X(_3687_));
 sky130_fd_sc_hd__nand2_1 _4592_ (.A(_1100_),
    .B(_3687_),
    .Y(_3688_));
 sky130_fd_sc_hd__mux2_1 _4593_ (.A0(_3675_),
    .A1(_3688_),
    .S(_1012_),
    .X(_3689_));
 sky130_fd_sc_hd__mux2_1 _4594_ (.A0(_3653_),
    .A1(_3689_),
    .S(_0957_),
    .X(_3690_));
 sky130_fd_sc_hd__mux2_1 _4595_ (.A0(_3091_),
    .A1(_3690_),
    .S(_0913_),
    .X(_3691_));
 sky130_fd_sc_hd__a21oi_1 _4596_ (.A1(_2024_),
    .A2(_2167_),
    .B1(_1672_),
    .Y(_3692_));
 sky130_fd_sc_hd__a21oi_1 _4597_ (.A1(_1441_),
    .A2(_3691_),
    .B1(_3692_),
    .Y(_3693_));
 sky130_fd_sc_hd__mux2_1 _4598_ (.A0(net58),
    .A1(_3693_),
    .S(_0814_),
    .X(_3694_));
 sky130_fd_sc_hd__inv_2 _4599_ (.A(_3694_),
    .Y(_3695_));
 sky130_fd_sc_hd__mux2_1 _4600_ (.A0(net26),
    .A1(_3693_),
    .S(_0858_),
    .X(_3696_));
 sky130_fd_sc_hd__or2_1 _4601_ (.A(_3695_),
    .B(_3696_),
    .X(_3697_));
 sky130_fd_sc_hd__nand2_1 _4602_ (.A(_1012_),
    .B(_1573_),
    .Y(_3698_));
 sky130_fd_sc_hd__o211a_1 _4603_ (.A1(_1012_),
    .A2(_1540_),
    .B1(_3698_),
    .C1(_0957_),
    .X(_3699_));
 sky130_fd_sc_hd__a21o_1 _4604_ (.A1(_0968_),
    .A2(_3643_),
    .B1(_3699_),
    .X(_3700_));
 sky130_fd_sc_hd__mux2_1 _4605_ (.A0(_3355_),
    .A1(_3700_),
    .S(_0913_),
    .X(_3701_));
 sky130_fd_sc_hd__o22a_1 _4606_ (.A1(_1672_),
    .A2(_2266_),
    .B1(_3701_),
    .B2(_1430_),
    .X(_3702_));
 sky130_fd_sc_hd__mux2_1 _4607_ (.A0(net55),
    .A1(_3702_),
    .S(_0814_),
    .X(_3703_));
 sky130_fd_sc_hd__or2_1 _4608_ (.A(_0869_),
    .B(_3702_),
    .X(_3704_));
 sky130_fd_sc_hd__o21ai_1 _4609_ (.A1(net23),
    .A2(_0858_),
    .B1(_3704_),
    .Y(_3705_));
 sky130_fd_sc_hd__inv_2 _4610_ (.A(_3705_),
    .Y(_3706_));
 sky130_fd_sc_hd__a2bb2o_1 _4611_ (.A1_N(_3705_),
    .A2_N(_3703_),
    .B1(_3696_),
    .B2(_3695_),
    .X(_3707_));
 sky130_fd_sc_hd__nor2_1 _4612_ (.A(_1012_),
    .B(_3688_),
    .Y(_3708_));
 sky130_fd_sc_hd__mux4_1 _4613_ (.A0(net44),
    .A1(net12),
    .A2(net55),
    .A3(net23),
    .S0(_1144_),
    .S1(_0649_),
    .X(_3709_));
 sky130_fd_sc_hd__a31o_1 _4614_ (.A1(_1012_),
    .A2(_1100_),
    .A3(_3709_),
    .B1(_0968_),
    .X(_3710_));
 sky130_fd_sc_hd__o221a_1 _4615_ (.A1(_0957_),
    .A2(_3676_),
    .B1(_3708_),
    .B2(_3710_),
    .C1(_0913_),
    .X(_3711_));
 sky130_fd_sc_hd__a211o_1 _4616_ (.A1(_0924_),
    .A2(_3457_),
    .B1(_3711_),
    .C1(_1430_),
    .X(_3712_));
 sky130_fd_sc_hd__a21o_1 _4617_ (.A1(_2024_),
    .A2(_2354_),
    .B1(_1672_),
    .X(_3713_));
 sky130_fd_sc_hd__and2_1 _4618_ (.A(_3712_),
    .B(_3713_),
    .X(_3714_));
 sky130_fd_sc_hd__mux2_1 _4619_ (.A0(net44),
    .A1(_3714_),
    .S(_0814_),
    .X(_3715_));
 sky130_fd_sc_hd__or2_1 _4620_ (.A(_0869_),
    .B(_3714_),
    .X(_3716_));
 sky130_fd_sc_hd__o21ai_2 _4621_ (.A1(net12),
    .A2(_0858_),
    .B1(_3716_),
    .Y(_3717_));
 sky130_fd_sc_hd__inv_2 _4622_ (.A(_3717_),
    .Y(_3718_));
 sky130_fd_sc_hd__a22o_1 _4623_ (.A1(_3703_),
    .A2(_3705_),
    .B1(_3715_),
    .B2(_3717_),
    .X(_3719_));
 sky130_fd_sc_hd__nand2b_1 _4624_ (.A_N(_2068_),
    .B(_2079_),
    .Y(_3720_));
 sky130_fd_sc_hd__o21a_1 _4625_ (.A1(_3715_),
    .A2(_3717_),
    .B1(_3720_),
    .X(_3721_));
 sky130_fd_sc_hd__o21ai_1 _4626_ (.A1(_3715_),
    .A2(_3717_),
    .B1(_3720_),
    .Y(_3722_));
 sky130_fd_sc_hd__o21bai_1 _4627_ (.A1(_3719_),
    .A2(_3721_),
    .B1_N(_3707_),
    .Y(_3723_));
 sky130_fd_sc_hd__a21oi_1 _4628_ (.A1(_3697_),
    .A2(_3723_),
    .B1(_3686_),
    .Y(_3724_));
 sky130_fd_sc_hd__nor2_1 _4629_ (.A(_3658_),
    .B(_3660_),
    .Y(_3725_));
 sky130_fd_sc_hd__a2bb2o_1 _4630_ (.A1_N(_3647_),
    .A2_N(_3649_),
    .B1(_3681_),
    .B2(_3683_),
    .X(_3726_));
 sky130_fd_sc_hd__a21oi_1 _4631_ (.A1(_3663_),
    .A2(_3726_),
    .B1(_3725_),
    .Y(_3727_));
 sky130_fd_sc_hd__xor2_1 _4632_ (.A(_3563_),
    .B(_3573_),
    .X(_3728_));
 sky130_fd_sc_hd__or4_1 _4633_ (.A(_3025_),
    .B(_3419_),
    .C(_3534_),
    .D(_3728_),
    .X(_3729_));
 sky130_fd_sc_hd__o2111a_1 _4634_ (.A1(_2992_),
    .A2(_3014_),
    .B1(_3524_),
    .C1(_3603_),
    .D1(_2926_),
    .X(_3730_));
 sky130_fd_sc_hd__nand2_1 _4635_ (.A(_3613_),
    .B(_3730_),
    .Y(_3731_));
 sky130_fd_sc_hd__nor2_1 _4636_ (.A(_3729_),
    .B(_3731_),
    .Y(_3732_));
 sky130_fd_sc_hd__o211a_1 _4637_ (.A1(_3685_),
    .A2(_3724_),
    .B1(_3727_),
    .C1(_3732_),
    .X(_3733_));
 sky130_fd_sc_hd__a21o_1 _4638_ (.A1(_2926_),
    .A2(_3641_),
    .B1(_3733_),
    .X(_3734_));
 sky130_fd_sc_hd__and2_1 _4639_ (.A(_2783_),
    .B(_3734_),
    .X(_3735_));
 sky130_fd_sc_hd__and3b_1 _4640_ (.A_N(_2299_),
    .B(_2288_),
    .C(_2211_),
    .X(_3736_));
 sky130_fd_sc_hd__a211o_1 _4641_ (.A1(_2420_),
    .A2(_2695_),
    .B1(_3736_),
    .C1(_2574_),
    .X(_3737_));
 sky130_fd_sc_hd__a21o_1 _4642_ (.A1(_2706_),
    .A2(_3737_),
    .B1(_2563_),
    .X(_3738_));
 sky130_fd_sc_hd__a221o_1 _4643_ (.A1(_0803_),
    .A2(_2728_),
    .B1(_2739_),
    .B2(_3738_),
    .C1(_3735_),
    .X(_3739_));
 sky130_fd_sc_hd__nand2b_1 _4644_ (.A_N(_2079_),
    .B(_2068_),
    .Y(_3740_));
 sky130_fd_sc_hd__or4_1 _4645_ (.A(_3707_),
    .B(_3719_),
    .C(_3722_),
    .D(_3726_),
    .X(_3741_));
 sky130_fd_sc_hd__or4b_1 _4646_ (.A(_2794_),
    .B(_3685_),
    .C(_3725_),
    .D_N(_3740_),
    .X(_3742_));
 sky130_fd_sc_hd__or4b_1 _4647_ (.A(_3686_),
    .B(_3741_),
    .C(_3742_),
    .D_N(_3697_),
    .X(_3743_));
 sky130_fd_sc_hd__o31a_4 _4648_ (.A1(_3729_),
    .A2(_3731_),
    .A3(_3743_),
    .B1(_3739_),
    .X(_3744_));
 sky130_fd_sc_hd__xor2_4 _4649_ (.A(net25),
    .B(net57),
    .X(_3745_));
 sky130_fd_sc_hd__xnor2_4 _4650_ (.A(net25),
    .B(net57),
    .Y(_3746_));
 sky130_fd_sc_hd__mux2_1 _4651_ (.A0(_2068_),
    .A1(_2079_),
    .S(_3744_),
    .X(_3747_));
 sky130_fd_sc_hd__nand2_1 _4652_ (.A(_3745_),
    .B(_3747_),
    .Y(_3748_));
 sky130_fd_sc_hd__mux2_1 _4653_ (.A0(_3715_),
    .A1(_3718_),
    .S(_3744_),
    .X(_3749_));
 sky130_fd_sc_hd__xnor2_1 _4654_ (.A(_3748_),
    .B(_3749_),
    .Y(_3750_));
 sky130_fd_sc_hd__mux2_1 _4655_ (.A0(_3718_),
    .A1(_3715_),
    .S(_3744_),
    .X(_3751_));
 sky130_fd_sc_hd__xnor2_1 _4656_ (.A(_3750_),
    .B(_3751_),
    .Y(_3752_));
 sky130_fd_sc_hd__xnor2_2 _4657_ (.A(_2090_),
    .B(_3752_),
    .Y(_3753_));
 sky130_fd_sc_hd__or2_1 _4658_ (.A(_1430_),
    .B(_3656_),
    .X(_3754_));
 sky130_fd_sc_hd__o21a_1 _4659_ (.A1(_3747_),
    .A2(_3749_),
    .B1(_3745_),
    .X(_3755_));
 sky130_fd_sc_hd__mux2_1 _4660_ (.A0(_3703_),
    .A1(_3706_),
    .S(_3744_),
    .X(_3756_));
 sky130_fd_sc_hd__nor2_1 _4661_ (.A(_3755_),
    .B(_3756_),
    .Y(_3757_));
 sky130_fd_sc_hd__inv_2 _4662_ (.A(_3757_),
    .Y(_3758_));
 sky130_fd_sc_hd__mux2_1 _4663_ (.A0(_3694_),
    .A1(_3696_),
    .S(_3744_),
    .X(_3759_));
 sky130_fd_sc_hd__mux2_1 _4664_ (.A0(_3669_),
    .A1(_3671_),
    .S(_3744_),
    .X(_3760_));
 sky130_fd_sc_hd__mux2_1 _4665_ (.A0(_3681_),
    .A1(_3684_),
    .S(_3744_),
    .X(_3761_));
 sky130_fd_sc_hd__or4b_1 _4666_ (.A(_3758_),
    .B(_3759_),
    .C(_3760_),
    .D_N(_3761_),
    .X(_3762_));
 sky130_fd_sc_hd__mux2_1 _4667_ (.A0(_3647_),
    .A1(_3648_),
    .S(_3744_),
    .X(_3763_));
 sky130_fd_sc_hd__mux2_1 _4668_ (.A0(_3658_),
    .A1(_3661_),
    .S(_3744_),
    .X(_3764_));
 sky130_fd_sc_hd__mux2_1 _4669_ (.A0(_3563_),
    .A1(_3573_),
    .S(_3744_),
    .X(_3765_));
 sky130_fd_sc_hd__or4_1 _4670_ (.A(_3762_),
    .B(_3763_),
    .C(_3764_),
    .D(_3765_),
    .X(_3766_));
 sky130_fd_sc_hd__mux2_1 _4671_ (.A0(_3505_),
    .A1(_3515_),
    .S(_3744_),
    .X(_3767_));
 sky130_fd_sc_hd__or2_1 _4672_ (.A(_3766_),
    .B(_3767_),
    .X(_3768_));
 sky130_fd_sc_hd__mux2_1 _4673_ (.A0(_3386_),
    .A1(_3408_),
    .S(_3744_),
    .X(_3769_));
 sky130_fd_sc_hd__or2_1 _4674_ (.A(_3768_),
    .B(_3769_),
    .X(_3770_));
 sky130_fd_sc_hd__mux2_1 _4675_ (.A0(_3124_),
    .A1(_3146_),
    .S(_3744_),
    .X(_3771_));
 sky130_fd_sc_hd__nor2_1 _4676_ (.A(_3770_),
    .B(_3771_),
    .Y(_3772_));
 sky130_fd_sc_hd__inv_2 _4677_ (.A(_3772_),
    .Y(_3773_));
 sky130_fd_sc_hd__mux2_1 _4678_ (.A0(_3212_),
    .A1(_3223_),
    .S(_3744_),
    .X(_3774_));
 sky130_fd_sc_hd__mux2_1 _4679_ (.A0(_3311_),
    .A1(_3322_),
    .S(_3744_),
    .X(_3775_));
 sky130_fd_sc_hd__or3_1 _4680_ (.A(_3773_),
    .B(_3774_),
    .C(_3775_),
    .X(_3776_));
 sky130_fd_sc_hd__mux2_1 _4681_ (.A0(_2992_),
    .A1(_3003_),
    .S(_3744_),
    .X(_3777_));
 sky130_fd_sc_hd__nor2_1 _4682_ (.A(_3776_),
    .B(_3777_),
    .Y(_3778_));
 sky130_fd_sc_hd__mux2_1 _4683_ (.A0(_2904_),
    .A1(_2915_),
    .S(_3744_),
    .X(_3779_));
 sky130_fd_sc_hd__or3_1 _4684_ (.A(_3776_),
    .B(_3777_),
    .C(_3779_),
    .X(_3780_));
 sky130_fd_sc_hd__mux2_1 _4685_ (.A0(_2662_),
    .A1(_2673_),
    .S(_3744_),
    .X(_3781_));
 sky130_fd_sc_hd__mux2_1 _4686_ (.A0(_2376_),
    .A1(_2387_),
    .S(_3744_),
    .X(_3782_));
 sky130_fd_sc_hd__mux2_1 _4687_ (.A0(_2288_),
    .A1(_2299_),
    .S(_3744_),
    .X(_3783_));
 sky130_fd_sc_hd__or4_1 _4688_ (.A(_3780_),
    .B(_3781_),
    .C(_3782_),
    .D(_3783_),
    .X(_3784_));
 sky130_fd_sc_hd__mux2_1 _4689_ (.A0(_2189_),
    .A1(_2200_),
    .S(_3744_),
    .X(_3785_));
 sky130_fd_sc_hd__mux2_1 _4690_ (.A0(_2530_),
    .A1(_2541_),
    .S(_3744_),
    .X(_3786_));
 sky130_fd_sc_hd__mux2_1 _4691_ (.A0(_2464_),
    .A1(_2475_),
    .S(_3744_),
    .X(_3787_));
 sky130_fd_sc_hd__mux2_1 _4692_ (.A0(_2717_),
    .A1(_2618_),
    .S(_3744_),
    .X(_3788_));
 sky130_fd_sc_hd__nor2_1 _4693_ (.A(_3746_),
    .B(_3757_),
    .Y(_3789_));
 sky130_fd_sc_hd__a21oi_1 _4694_ (.A1(_3745_),
    .A2(_3759_),
    .B1(_3789_),
    .Y(_3790_));
 sky130_fd_sc_hd__a21boi_1 _4695_ (.A1(_3745_),
    .A2(_3760_),
    .B1_N(_3790_),
    .Y(_3791_));
 sky130_fd_sc_hd__and2_1 _4696_ (.A(_3745_),
    .B(_3762_),
    .X(_3792_));
 sky130_fd_sc_hd__o21a_1 _4697_ (.A1(_3762_),
    .A2(_3763_),
    .B1(_3745_),
    .X(_3793_));
 sky130_fd_sc_hd__a21o_1 _4698_ (.A1(_3745_),
    .A2(_3764_),
    .B1(_3793_),
    .X(_3794_));
 sky130_fd_sc_hd__nand2_1 _4699_ (.A(_3745_),
    .B(_3766_),
    .Y(_3795_));
 sky130_fd_sc_hd__and2_1 _4700_ (.A(_3745_),
    .B(_3768_),
    .X(_3796_));
 sky130_fd_sc_hd__and2_1 _4701_ (.A(_3745_),
    .B(_3770_),
    .X(_3797_));
 sky130_fd_sc_hd__or2_1 _4702_ (.A(_3746_),
    .B(_3772_),
    .X(_3798_));
 sky130_fd_sc_hd__o21a_1 _4703_ (.A1(_3773_),
    .A2(_3774_),
    .B1(_3745_),
    .X(_3799_));
 sky130_fd_sc_hd__and2_1 _4704_ (.A(_3745_),
    .B(_3776_),
    .X(_3800_));
 sky130_fd_sc_hd__nor2_1 _4705_ (.A(_3746_),
    .B(_3778_),
    .Y(_3801_));
 sky130_fd_sc_hd__and2_1 _4706_ (.A(_3745_),
    .B(_3780_),
    .X(_3802_));
 sky130_fd_sc_hd__o21a_1 _4707_ (.A1(_3780_),
    .A2(_3781_),
    .B1(_3745_),
    .X(_3803_));
 sky130_fd_sc_hd__a21o_1 _4708_ (.A1(_3745_),
    .A2(_3782_),
    .B1(_3803_),
    .X(_3804_));
 sky130_fd_sc_hd__and2_1 _4709_ (.A(_3745_),
    .B(_3784_),
    .X(_3805_));
 sky130_fd_sc_hd__o21a_1 _4710_ (.A1(_3784_),
    .A2(_3785_),
    .B1(_3745_),
    .X(_3806_));
 sky130_fd_sc_hd__a21oi_1 _4711_ (.A1(_3745_),
    .A2(_3786_),
    .B1(_3806_),
    .Y(_3807_));
 sky130_fd_sc_hd__a21bo_1 _4712_ (.A1(_3745_),
    .A2(_3787_),
    .B1_N(_3807_),
    .X(_3808_));
 sky130_fd_sc_hd__a21oi_1 _4713_ (.A1(_3745_),
    .A2(_3788_),
    .B1(_3808_),
    .Y(_3809_));
 sky130_fd_sc_hd__xor2_1 _4714_ (.A(_3754_),
    .B(_3809_),
    .X(_3810_));
 sky130_fd_sc_hd__o21a_1 _4715_ (.A1(net98),
    .A2(_1760_),
    .B1(_3810_),
    .X(_3811_));
 sky130_fd_sc_hd__and3b_1 _4716_ (.A_N(_3810_),
    .B(_1771_),
    .C(_0803_),
    .X(_3812_));
 sky130_fd_sc_hd__nor2_1 _4717_ (.A(_3811_),
    .B(_3812_),
    .Y(_3813_));
 sky130_fd_sc_hd__xnor2_1 _4718_ (.A(_3788_),
    .B(_3808_),
    .Y(_3814_));
 sky130_fd_sc_hd__mux2_1 _4719_ (.A0(_2618_),
    .A1(_2717_),
    .S(_3744_),
    .X(_3815_));
 sky130_fd_sc_hd__nand2b_1 _4720_ (.A_N(_3814_),
    .B(_3815_),
    .Y(_3816_));
 sky130_fd_sc_hd__xor2_2 _4721_ (.A(_3814_),
    .B(_3815_),
    .X(_3817_));
 sky130_fd_sc_hd__xnor2_1 _4722_ (.A(_3787_),
    .B(_3807_),
    .Y(_3818_));
 sky130_fd_sc_hd__mux2_1 _4723_ (.A0(_2475_),
    .A1(_2464_),
    .S(_3744_),
    .X(_3819_));
 sky130_fd_sc_hd__xnor2_1 _4724_ (.A(_3818_),
    .B(_3819_),
    .Y(_3820_));
 sky130_fd_sc_hd__xor2_1 _4725_ (.A(_3786_),
    .B(_3806_),
    .X(_3821_));
 sky130_fd_sc_hd__mux2_1 _4726_ (.A0(_2541_),
    .A1(_2530_),
    .S(_3744_),
    .X(_3822_));
 sky130_fd_sc_hd__nand2_1 _4727_ (.A(_3821_),
    .B(_3822_),
    .Y(_3823_));
 sky130_fd_sc_hd__or2_1 _4728_ (.A(_3821_),
    .B(_3822_),
    .X(_3824_));
 sky130_fd_sc_hd__and2_1 _4729_ (.A(_3823_),
    .B(_3824_),
    .X(_3825_));
 sky130_fd_sc_hd__xor2_1 _4730_ (.A(_3785_),
    .B(_3805_),
    .X(_3826_));
 sky130_fd_sc_hd__mux2_1 _4731_ (.A0(_2200_),
    .A1(_2189_),
    .S(_3744_),
    .X(_3827_));
 sky130_fd_sc_hd__and2_1 _4732_ (.A(_3826_),
    .B(_3827_),
    .X(_3828_));
 sky130_fd_sc_hd__nor2_1 _4733_ (.A(_3826_),
    .B(_3827_),
    .Y(_3829_));
 sky130_fd_sc_hd__or2_1 _4734_ (.A(_3828_),
    .B(_3829_),
    .X(_3830_));
 sky130_fd_sc_hd__xor2_1 _4735_ (.A(_3783_),
    .B(_3804_),
    .X(_3831_));
 sky130_fd_sc_hd__mux2_1 _4736_ (.A0(_2299_),
    .A1(_2288_),
    .S(_3744_),
    .X(_3832_));
 sky130_fd_sc_hd__xnor2_1 _4737_ (.A(_3831_),
    .B(_3832_),
    .Y(_3833_));
 sky130_fd_sc_hd__xor2_1 _4738_ (.A(_3782_),
    .B(_3803_),
    .X(_3834_));
 sky130_fd_sc_hd__mux2_1 _4739_ (.A0(_2387_),
    .A1(_2376_),
    .S(_3744_),
    .X(_3835_));
 sky130_fd_sc_hd__nand2_1 _4740_ (.A(_3834_),
    .B(_3835_),
    .Y(_3836_));
 sky130_fd_sc_hd__or2_1 _4741_ (.A(_3834_),
    .B(_3835_),
    .X(_3837_));
 sky130_fd_sc_hd__and2_1 _4742_ (.A(_3836_),
    .B(_3837_),
    .X(_3838_));
 sky130_fd_sc_hd__xnor2_1 _4743_ (.A(_3781_),
    .B(_3802_),
    .Y(_3839_));
 sky130_fd_sc_hd__mux2_1 _4744_ (.A0(_2673_),
    .A1(_2662_),
    .S(_3744_),
    .X(_3840_));
 sky130_fd_sc_hd__and2b_1 _4745_ (.A_N(_3839_),
    .B(_3840_),
    .X(_3841_));
 sky130_fd_sc_hd__xnor2_1 _4746_ (.A(_3839_),
    .B(_3840_),
    .Y(_3842_));
 sky130_fd_sc_hd__xnor2_1 _4747_ (.A(_3779_),
    .B(_3801_),
    .Y(_3843_));
 sky130_fd_sc_hd__mux2_1 _4748_ (.A0(_2915_),
    .A1(_2904_),
    .S(_3744_),
    .X(_3844_));
 sky130_fd_sc_hd__and2b_1 _4749_ (.A_N(_3843_),
    .B(_3844_),
    .X(_3845_));
 sky130_fd_sc_hd__xor2_1 _4750_ (.A(_3843_),
    .B(_3844_),
    .X(_3846_));
 sky130_fd_sc_hd__xnor2_1 _4751_ (.A(_3777_),
    .B(_3800_),
    .Y(_3847_));
 sky130_fd_sc_hd__mux2_1 _4752_ (.A0(_3003_),
    .A1(_2992_),
    .S(_3744_),
    .X(_3848_));
 sky130_fd_sc_hd__nand2b_1 _4753_ (.A_N(_3847_),
    .B(_3848_),
    .Y(_3849_));
 sky130_fd_sc_hd__xor2_1 _4754_ (.A(_3847_),
    .B(_3848_),
    .X(_3850_));
 sky130_fd_sc_hd__xor2_1 _4755_ (.A(_3775_),
    .B(_3799_),
    .X(_3851_));
 sky130_fd_sc_hd__mux2_1 _4756_ (.A0(_3322_),
    .A1(_3311_),
    .S(_3744_),
    .X(_3852_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(_3851_),
    .B(_3852_),
    .Y(_3853_));
 sky130_fd_sc_hd__or2_1 _4758_ (.A(_3851_),
    .B(_3852_),
    .X(_3854_));
 sky130_fd_sc_hd__and2_1 _4759_ (.A(_3853_),
    .B(_3854_),
    .X(_3855_));
 sky130_fd_sc_hd__xnor2_1 _4760_ (.A(_3774_),
    .B(_3798_),
    .Y(_3856_));
 sky130_fd_sc_hd__mux2_1 _4761_ (.A0(_3223_),
    .A1(_3212_),
    .S(_3744_),
    .X(_3857_));
 sky130_fd_sc_hd__and2_1 _4762_ (.A(_3856_),
    .B(_3857_),
    .X(_3858_));
 sky130_fd_sc_hd__nor2_1 _4763_ (.A(_3856_),
    .B(_3857_),
    .Y(_3859_));
 sky130_fd_sc_hd__or2_1 _4764_ (.A(_3858_),
    .B(_3859_),
    .X(_3860_));
 sky130_fd_sc_hd__xnor2_1 _4765_ (.A(_3771_),
    .B(_3797_),
    .Y(_3861_));
 sky130_fd_sc_hd__inv_2 _4766_ (.A(_3861_),
    .Y(_3862_));
 sky130_fd_sc_hd__mux2_1 _4767_ (.A0(_3146_),
    .A1(_3124_),
    .S(_3744_),
    .X(_3863_));
 sky130_fd_sc_hd__xnor2_1 _4768_ (.A(_3861_),
    .B(_3863_),
    .Y(_3864_));
 sky130_fd_sc_hd__xor2_1 _4769_ (.A(_3769_),
    .B(_3796_),
    .X(_3865_));
 sky130_fd_sc_hd__mux2_1 _4770_ (.A0(_3408_),
    .A1(_3386_),
    .S(_3744_),
    .X(_3866_));
 sky130_fd_sc_hd__and2_1 _4771_ (.A(_3865_),
    .B(_3866_),
    .X(_3867_));
 sky130_fd_sc_hd__nor2_1 _4772_ (.A(_3865_),
    .B(_3866_),
    .Y(_3868_));
 sky130_fd_sc_hd__or2_1 _4773_ (.A(_3867_),
    .B(_3868_),
    .X(_3869_));
 sky130_fd_sc_hd__xnor2_1 _4774_ (.A(_3767_),
    .B(_3795_),
    .Y(_3870_));
 sky130_fd_sc_hd__mux2_1 _4775_ (.A0(_3515_),
    .A1(_3505_),
    .S(_3744_),
    .X(_3871_));
 sky130_fd_sc_hd__xnor2_1 _4776_ (.A(_3870_),
    .B(_3871_),
    .Y(_3872_));
 sky130_fd_sc_hd__xnor2_2 _4777_ (.A(_3765_),
    .B(_3794_),
    .Y(_3873_));
 sky130_fd_sc_hd__mux2_1 _4778_ (.A0(_3573_),
    .A1(_3563_),
    .S(_3744_),
    .X(_3874_));
 sky130_fd_sc_hd__nand2b_1 _4779_ (.A_N(_3873_),
    .B(_3874_),
    .Y(_3875_));
 sky130_fd_sc_hd__xor2_2 _4780_ (.A(_3873_),
    .B(_3874_),
    .X(_3876_));
 sky130_fd_sc_hd__xnor2_1 _4781_ (.A(_3764_),
    .B(_3793_),
    .Y(_3877_));
 sky130_fd_sc_hd__mux2_1 _4782_ (.A0(_3661_),
    .A1(_3658_),
    .S(_3744_),
    .X(_3878_));
 sky130_fd_sc_hd__nand2b_1 _4783_ (.A_N(_3877_),
    .B(_3878_),
    .Y(_3879_));
 sky130_fd_sc_hd__xnor2_1 _4784_ (.A(_3877_),
    .B(_3878_),
    .Y(_3880_));
 sky130_fd_sc_hd__xnor2_1 _4785_ (.A(_3763_),
    .B(_3792_),
    .Y(_3881_));
 sky130_fd_sc_hd__mux2_1 _4786_ (.A0(_3648_),
    .A1(_3647_),
    .S(_3744_),
    .X(_3882_));
 sky130_fd_sc_hd__and2b_1 _4787_ (.A_N(_3881_),
    .B(_3882_),
    .X(_3883_));
 sky130_fd_sc_hd__xor2_1 _4788_ (.A(_3881_),
    .B(_3882_),
    .X(_3884_));
 sky130_fd_sc_hd__xor2_1 _4789_ (.A(_3761_),
    .B(_3791_),
    .X(_3885_));
 sky130_fd_sc_hd__mux2_1 _4790_ (.A0(_3683_),
    .A1(_3682_),
    .S(_3744_),
    .X(_3886_));
 sky130_fd_sc_hd__xnor2_1 _4791_ (.A(_3885_),
    .B(_3886_),
    .Y(_3887_));
 sky130_fd_sc_hd__xor2_1 _4792_ (.A(_3760_),
    .B(_3790_),
    .X(_3888_));
 sky130_fd_sc_hd__mux2_1 _4793_ (.A0(_3671_),
    .A1(_3669_),
    .S(_3744_),
    .X(_3889_));
 sky130_fd_sc_hd__nand2b_1 _4794_ (.A_N(_3888_),
    .B(_3889_),
    .Y(_3890_));
 sky130_fd_sc_hd__xor2_1 _4795_ (.A(_3888_),
    .B(_3889_),
    .X(_3891_));
 sky130_fd_sc_hd__xnor2_1 _4796_ (.A(_3759_),
    .B(_3789_),
    .Y(_3892_));
 sky130_fd_sc_hd__mux2_1 _4797_ (.A0(_3696_),
    .A1(_3694_),
    .S(_3744_),
    .X(_3893_));
 sky130_fd_sc_hd__nand2b_1 _4798_ (.A_N(_3892_),
    .B(_3893_),
    .Y(_3894_));
 sky130_fd_sc_hd__nand2b_1 _4799_ (.A_N(_3893_),
    .B(_3892_),
    .Y(_3895_));
 sky130_fd_sc_hd__nand2_1 _4800_ (.A(_3894_),
    .B(_3895_),
    .Y(_3896_));
 sky130_fd_sc_hd__xor2_1 _4801_ (.A(_3755_),
    .B(_3756_),
    .X(_3897_));
 sky130_fd_sc_hd__mux2_1 _4802_ (.A0(_3706_),
    .A1(_3703_),
    .S(_3744_),
    .X(_3898_));
 sky130_fd_sc_hd__nand2_1 _4803_ (.A(_3897_),
    .B(_3898_),
    .Y(_3899_));
 sky130_fd_sc_hd__a2bb2o_1 _4804_ (.A1_N(_2090_),
    .A2_N(_3752_),
    .B1(_3751_),
    .B2(_3750_),
    .X(_3900_));
 sky130_fd_sc_hd__or2_1 _4805_ (.A(_3897_),
    .B(_3898_),
    .X(_3901_));
 sky130_fd_sc_hd__nand2_1 _4806_ (.A(_3899_),
    .B(_3901_),
    .Y(_3902_));
 sky130_fd_sc_hd__nand2b_1 _4807_ (.A_N(_3902_),
    .B(_3900_),
    .Y(_3903_));
 sky130_fd_sc_hd__a21o_1 _4808_ (.A1(_3899_),
    .A2(_3903_),
    .B1(_3896_),
    .X(_3904_));
 sky130_fd_sc_hd__a21o_1 _4809_ (.A1(_3894_),
    .A2(_3904_),
    .B1(_3891_),
    .X(_3905_));
 sky130_fd_sc_hd__a21oi_1 _4810_ (.A1(_3890_),
    .A2(_3905_),
    .B1(_3887_),
    .Y(_3906_));
 sky130_fd_sc_hd__a21o_1 _4811_ (.A1(_3885_),
    .A2(_3886_),
    .B1(_3906_),
    .X(_3907_));
 sky130_fd_sc_hd__and2b_1 _4812_ (.A_N(_3884_),
    .B(_3907_),
    .X(_3908_));
 sky130_fd_sc_hd__o21ai_1 _4813_ (.A1(_3883_),
    .A2(_3908_),
    .B1(_3880_),
    .Y(_3909_));
 sky130_fd_sc_hd__nand2_1 _4814_ (.A(_3879_),
    .B(_3909_),
    .Y(_3910_));
 sky130_fd_sc_hd__a21o_1 _4815_ (.A1(_3879_),
    .A2(_3909_),
    .B1(_3876_),
    .X(_3911_));
 sky130_fd_sc_hd__a21oi_1 _4816_ (.A1(_3875_),
    .A2(_3911_),
    .B1(_3872_),
    .Y(_3912_));
 sky130_fd_sc_hd__a21o_1 _4817_ (.A1(_3870_),
    .A2(_3871_),
    .B1(_3912_),
    .X(_3913_));
 sky130_fd_sc_hd__and2b_1 _4818_ (.A_N(_3869_),
    .B(_3913_),
    .X(_3914_));
 sky130_fd_sc_hd__o21ai_1 _4819_ (.A1(_3867_),
    .A2(_3914_),
    .B1(_3864_),
    .Y(_3915_));
 sky130_fd_sc_hd__a21boi_2 _4820_ (.A1(_3862_),
    .A2(_3863_),
    .B1_N(_3915_),
    .Y(_3916_));
 sky130_fd_sc_hd__nor2_1 _4821_ (.A(_3860_),
    .B(_3916_),
    .Y(_3917_));
 sky130_fd_sc_hd__o21ai_1 _4822_ (.A1(_3858_),
    .A2(_3917_),
    .B1(_3855_),
    .Y(_3918_));
 sky130_fd_sc_hd__a21o_1 _4823_ (.A1(_3853_),
    .A2(_3918_),
    .B1(_3850_),
    .X(_3919_));
 sky130_fd_sc_hd__a21oi_1 _4824_ (.A1(_3849_),
    .A2(_3919_),
    .B1(_3846_),
    .Y(_3920_));
 sky130_fd_sc_hd__o21a_1 _4825_ (.A1(_3845_),
    .A2(_3920_),
    .B1(_3842_),
    .X(_3921_));
 sky130_fd_sc_hd__o21ai_1 _4826_ (.A1(_3841_),
    .A2(_3921_),
    .B1(_3838_),
    .Y(_3922_));
 sky130_fd_sc_hd__a21oi_1 _4827_ (.A1(_3836_),
    .A2(_3922_),
    .B1(_3833_),
    .Y(_3923_));
 sky130_fd_sc_hd__a21oi_1 _4828_ (.A1(_3831_),
    .A2(_3832_),
    .B1(_3923_),
    .Y(_3924_));
 sky130_fd_sc_hd__nor2_1 _4829_ (.A(_3830_),
    .B(_3924_),
    .Y(_3925_));
 sky130_fd_sc_hd__o21ai_1 _4830_ (.A1(_3828_),
    .A2(_3925_),
    .B1(_3825_),
    .Y(_3926_));
 sky130_fd_sc_hd__a21oi_1 _4831_ (.A1(_3823_),
    .A2(_3926_),
    .B1(_3820_),
    .Y(_3927_));
 sky130_fd_sc_hd__a21oi_2 _4832_ (.A1(_3818_),
    .A2(_3819_),
    .B1(_3927_),
    .Y(_3928_));
 sky130_fd_sc_hd__o21a_1 _4833_ (.A1(_3817_),
    .A2(_3928_),
    .B1(_3816_),
    .X(_3929_));
 sky130_fd_sc_hd__and2b_1 _4834_ (.A_N(_3929_),
    .B(_3813_),
    .X(_3930_));
 sky130_fd_sc_hd__a21o_1 _4835_ (.A1(_3754_),
    .A2(_3809_),
    .B1(_3746_),
    .X(_3931_));
 sky130_fd_sc_hd__o21a_4 _4836_ (.A1(_3811_),
    .A2(_3930_),
    .B1(_3931_),
    .X(_3932_));
 sky130_fd_sc_hd__clkinv_4 _4837_ (.A(_3932_),
    .Y(_3933_));
 sky130_fd_sc_hd__nand2_1 _4838_ (.A(_3720_),
    .B(_3740_),
    .Y(_3934_));
 sky130_fd_sc_hd__and2b_1 _4839_ (.A_N(_3813_),
    .B(_3929_),
    .X(_3935_));
 sky130_fd_sc_hd__nor2_2 _4840_ (.A(_3930_),
    .B(_3935_),
    .Y(_3936_));
 sky130_fd_sc_hd__or2_4 _4841_ (.A(_3930_),
    .B(_3935_),
    .X(_3937_));
 sky130_fd_sc_hd__nor2_4 _4842_ (.A(_3932_),
    .B(_3937_),
    .Y(_3938_));
 sky130_fd_sc_hd__or2_2 _4843_ (.A(_3932_),
    .B(_3937_),
    .X(_3939_));
 sky130_fd_sc_hd__o2bb2a_1 _4844_ (.A1_N(_3934_),
    .A2_N(_3938_),
    .B1(_3753_),
    .B2(_3933_),
    .X(_3940_));
 sky130_fd_sc_hd__or3_1 _4845_ (.A(_0308_),
    .B(_0451_),
    .C(_3746_),
    .X(_3941_));
 sky130_fd_sc_hd__o211a_1 _4846_ (.A1(_0462_),
    .A2(_3940_),
    .B1(_3941_),
    .C1(_1111_),
    .X(_3942_));
 sky130_fd_sc_hd__nor2_1 _4847_ (.A(net65),
    .B(_3942_),
    .Y(_3943_));
 sky130_fd_sc_hd__nand2_2 _4848_ (.A(_0297_),
    .B(_1771_),
    .Y(_3944_));
 sky130_fd_sc_hd__nand2_2 _4849_ (.A(_0396_),
    .B(_1727_),
    .Y(_3945_));
 sky130_fd_sc_hd__o221ai_2 _4850_ (.A1(_0451_),
    .A2(_3944_),
    .B1(_3945_),
    .B2(_0308_),
    .C1(_1111_),
    .Y(_3946_));
 sky130_fd_sc_hd__nor2_1 _4851_ (.A(_0176_),
    .B(_3946_),
    .Y(_3947_));
 sky130_fd_sc_hd__and3_1 _4852_ (.A(net21),
    .B(net53),
    .C(_0506_),
    .X(_3948_));
 sky130_fd_sc_hd__a21oi_1 _4853_ (.A1(net21),
    .A2(net53),
    .B1(_0506_),
    .Y(_3949_));
 sky130_fd_sc_hd__nor2_1 _4854_ (.A(_3948_),
    .B(_3949_),
    .Y(_3950_));
 sky130_fd_sc_hd__a21oi_1 _4855_ (.A1(net20),
    .A2(net52),
    .B1(_0825_),
    .Y(_3951_));
 sky130_fd_sc_hd__a21o_1 _4856_ (.A1(net20),
    .A2(net52),
    .B1(_0825_),
    .X(_3952_));
 sky130_fd_sc_hd__and3_1 _4857_ (.A(net20),
    .B(net52),
    .C(_0825_),
    .X(_3953_));
 sky130_fd_sc_hd__or2_1 _4858_ (.A(_3951_),
    .B(_3953_),
    .X(_3954_));
 sky130_fd_sc_hd__and3_1 _4859_ (.A(net18),
    .B(net50),
    .C(_0693_),
    .X(_3955_));
 sky130_fd_sc_hd__a21oi_1 _4860_ (.A1(net18),
    .A2(net50),
    .B1(_0693_),
    .Y(_3956_));
 sky130_fd_sc_hd__nor2_1 _4861_ (.A(_3955_),
    .B(_3956_),
    .Y(_3957_));
 sky130_fd_sc_hd__and3_1 _4862_ (.A(net17),
    .B(net49),
    .C(_0682_),
    .X(_3958_));
 sky130_fd_sc_hd__a21oi_1 _4863_ (.A1(net17),
    .A2(net49),
    .B1(_0682_),
    .Y(_3959_));
 sky130_fd_sc_hd__nor2_1 _4864_ (.A(_3958_),
    .B(_3959_),
    .Y(_3960_));
 sky130_fd_sc_hd__o21a_1 _4865_ (.A1(net16),
    .A2(net48),
    .B1(_0616_),
    .X(_3961_));
 sky130_fd_sc_hd__a21oi_1 _4866_ (.A1(_3960_),
    .A2(_3961_),
    .B1(_3958_),
    .Y(_3962_));
 sky130_fd_sc_hd__o21ba_1 _4867_ (.A1(_3956_),
    .A2(_3962_),
    .B1_N(_3955_),
    .X(_3963_));
 sky130_fd_sc_hd__and3_1 _4868_ (.A(net19),
    .B(net51),
    .C(_0572_),
    .X(_3964_));
 sky130_fd_sc_hd__a21oi_1 _4869_ (.A1(net19),
    .A2(net51),
    .B1(_0572_),
    .Y(_3965_));
 sky130_fd_sc_hd__or2_1 _4870_ (.A(_3964_),
    .B(_3965_),
    .X(_3966_));
 sky130_fd_sc_hd__nor2_1 _4871_ (.A(_3963_),
    .B(_3966_),
    .Y(_3967_));
 sky130_fd_sc_hd__o31ai_2 _4872_ (.A1(_3953_),
    .A2(_3964_),
    .A3(_3967_),
    .B1(_3952_),
    .Y(_3968_));
 sky130_fd_sc_hd__inv_2 _4873_ (.A(_3968_),
    .Y(_3969_));
 sky130_fd_sc_hd__xnor2_1 _4874_ (.A(_3950_),
    .B(_3968_),
    .Y(_3970_));
 sky130_fd_sc_hd__nor2_1 _4875_ (.A(net48),
    .B(_0616_),
    .Y(_3971_));
 sky130_fd_sc_hd__a21oi_1 _4876_ (.A1(_0121_),
    .A2(_3971_),
    .B1(_3961_),
    .Y(_3972_));
 sky130_fd_sc_hd__nand2_1 _4877_ (.A(net47),
    .B(_1716_),
    .Y(_3973_));
 sky130_fd_sc_hd__nand2_1 _4878_ (.A(net45),
    .B(_1716_),
    .Y(_3974_));
 sky130_fd_sc_hd__nand2_1 _4879_ (.A(net15),
    .B(net45),
    .Y(_3975_));
 sky130_fd_sc_hd__nand2_1 _4880_ (.A(net42),
    .B(_1716_),
    .Y(_3976_));
 sky130_fd_sc_hd__nand2_1 _4881_ (.A(net15),
    .B(net42),
    .Y(_3977_));
 sky130_fd_sc_hd__nand2_1 _4882_ (.A(net41),
    .B(_1716_),
    .Y(_3978_));
 sky130_fd_sc_hd__nand2_1 _4883_ (.A(net15),
    .B(net40),
    .Y(_3979_));
 sky130_fd_sc_hd__nand2_1 _4884_ (.A(net15),
    .B(net38),
    .Y(_3980_));
 sky130_fd_sc_hd__nand2_1 _4885_ (.A(net36),
    .B(_1716_),
    .Y(_3981_));
 sky130_fd_sc_hd__nand2_1 _4886_ (.A(net15),
    .B(net36),
    .Y(_3982_));
 sky130_fd_sc_hd__nor2_1 _4887_ (.A(_0055_),
    .B(_1727_),
    .Y(_3983_));
 sky130_fd_sc_hd__nand2_1 _4888_ (.A(net34),
    .B(_1716_),
    .Y(_3984_));
 sky130_fd_sc_hd__nand2_1 _4889_ (.A(net15),
    .B(net34),
    .Y(_3985_));
 sky130_fd_sc_hd__nand2_1 _4890_ (.A(net15),
    .B(net63),
    .Y(_3986_));
 sky130_fd_sc_hd__nand2_1 _4891_ (.A(net61),
    .B(_1716_),
    .Y(_3987_));
 sky130_fd_sc_hd__nand2_1 _4892_ (.A(net15),
    .B(net61),
    .Y(_3988_));
 sky130_fd_sc_hd__nand2_1 _4893_ (.A(net59),
    .B(_1716_),
    .Y(_3989_));
 sky130_fd_sc_hd__nand2_1 _4894_ (.A(net15),
    .B(net59),
    .Y(_3990_));
 sky130_fd_sc_hd__and2_1 _4895_ (.A(net55),
    .B(_1716_),
    .X(_3991_));
 sky130_fd_sc_hd__and3_1 _4896_ (.A(net44),
    .B(net33),
    .C(net15),
    .X(_3992_));
 sky130_fd_sc_hd__and2_1 _4897_ (.A(_1716_),
    .B(_3992_),
    .X(_3993_));
 sky130_fd_sc_hd__a22o_1 _4898_ (.A1(net44),
    .A2(net15),
    .B1(_1716_),
    .B2(net33),
    .X(_3994_));
 sky130_fd_sc_hd__and2_1 _4899_ (.A(net14),
    .B(_3992_),
    .X(_3995_));
 sky130_fd_sc_hd__a22o_1 _4900_ (.A1(net33),
    .A2(net15),
    .B1(net14),
    .B2(net44),
    .X(_3996_));
 sky130_fd_sc_hd__and4_1 _4901_ (.A(net44),
    .B(net33),
    .C(net14),
    .D(net13),
    .X(_3997_));
 sky130_fd_sc_hd__nand4_1 _4902_ (.A(net44),
    .B(net33),
    .C(net14),
    .D(net13),
    .Y(_3998_));
 sky130_fd_sc_hd__a22oi_2 _4903_ (.A1(net33),
    .A2(net14),
    .B1(net13),
    .B2(net44),
    .Y(_3999_));
 sky130_fd_sc_hd__a22o_1 _4904_ (.A1(net33),
    .A2(net13),
    .B1(net11),
    .B2(net44),
    .X(_4000_));
 sky130_fd_sc_hd__nand4_2 _4905_ (.A(net44),
    .B(net33),
    .C(net13),
    .D(net11),
    .Y(_4001_));
 sky130_fd_sc_hd__a22oi_1 _4906_ (.A1(net33),
    .A2(net11),
    .B1(net10),
    .B2(net44),
    .Y(_4002_));
 sky130_fd_sc_hd__nand4_2 _4907_ (.A(net44),
    .B(net33),
    .C(net11),
    .D(net10),
    .Y(_4003_));
 sky130_fd_sc_hd__a22oi_1 _4908_ (.A1(net33),
    .A2(net10),
    .B1(net9),
    .B2(net44),
    .Y(_4004_));
 sky130_fd_sc_hd__nand4_2 _4909_ (.A(net44),
    .B(net33),
    .C(net10),
    .D(net9),
    .Y(_4005_));
 sky130_fd_sc_hd__a22o_1 _4910_ (.A1(net33),
    .A2(net9),
    .B1(net8),
    .B2(net44),
    .X(_4006_));
 sky130_fd_sc_hd__and3_1 _4911_ (.A(net44),
    .B(net33),
    .C(net8),
    .X(_4007_));
 sky130_fd_sc_hd__and2_1 _4912_ (.A(net9),
    .B(_4007_),
    .X(_4008_));
 sky130_fd_sc_hd__a22o_1 _4913_ (.A1(net33),
    .A2(net8),
    .B1(net7),
    .B2(net44),
    .X(_4009_));
 sky130_fd_sc_hd__and3_1 _4914_ (.A(net44),
    .B(net33),
    .C(net7),
    .X(_4010_));
 sky130_fd_sc_hd__and2_1 _4915_ (.A(net8),
    .B(_4010_),
    .X(_4011_));
 sky130_fd_sc_hd__nand2_1 _4916_ (.A(net6),
    .B(_4010_),
    .Y(_4012_));
 sky130_fd_sc_hd__a22oi_2 _4917_ (.A1(net33),
    .A2(net7),
    .B1(net6),
    .B2(net44),
    .Y(_4013_));
 sky130_fd_sc_hd__nand4_2 _4918_ (.A(net44),
    .B(net33),
    .C(net6),
    .D(net5),
    .Y(_4014_));
 sky130_fd_sc_hd__a22o_1 _4919_ (.A1(net33),
    .A2(net6),
    .B1(net5),
    .B2(net44),
    .X(_4015_));
 sky130_fd_sc_hd__inv_2 _4920_ (.A(_4015_),
    .Y(_4016_));
 sky130_fd_sc_hd__and4_1 _4921_ (.A(net44),
    .B(net33),
    .C(net5),
    .D(net4),
    .X(_4017_));
 sky130_fd_sc_hd__inv_2 _4922_ (.A(_4017_),
    .Y(_4018_));
 sky130_fd_sc_hd__a22oi_2 _4923_ (.A1(net33),
    .A2(net5),
    .B1(net4),
    .B2(net44),
    .Y(_4019_));
 sky130_fd_sc_hd__nand4_2 _4924_ (.A(net44),
    .B(net33),
    .C(net4),
    .D(net3),
    .Y(_4020_));
 sky130_fd_sc_hd__a22o_1 _4925_ (.A1(net33),
    .A2(net4),
    .B1(net3),
    .B2(net44),
    .X(_4021_));
 sky130_fd_sc_hd__inv_2 _4926_ (.A(_4021_),
    .Y(_4022_));
 sky130_fd_sc_hd__a22oi_2 _4927_ (.A1(net33),
    .A2(net3),
    .B1(net2),
    .B2(net44),
    .Y(_4023_));
 sky130_fd_sc_hd__and4_1 _4928_ (.A(net44),
    .B(net33),
    .C(net3),
    .D(net2),
    .X(_4024_));
 sky130_fd_sc_hd__inv_2 _4929_ (.A(_4024_),
    .Y(_4025_));
 sky130_fd_sc_hd__a22o_1 _4930_ (.A1(net33),
    .A2(net2),
    .B1(net32),
    .B2(net44),
    .X(_4026_));
 sky130_fd_sc_hd__nand4_2 _4931_ (.A(net44),
    .B(net33),
    .C(net2),
    .D(net32),
    .Y(_4027_));
 sky130_fd_sc_hd__and4_1 _4932_ (.A(net44),
    .B(net33),
    .C(net32),
    .D(net31),
    .X(_4028_));
 sky130_fd_sc_hd__a22o_1 _4933_ (.A1(net33),
    .A2(net32),
    .B1(net31),
    .B2(net44),
    .X(_4029_));
 sky130_fd_sc_hd__and4_1 _4934_ (.A(net44),
    .B(net33),
    .C(net31),
    .D(net30),
    .X(_4030_));
 sky130_fd_sc_hd__nand4_1 _4935_ (.A(net44),
    .B(net33),
    .C(net31),
    .D(net30),
    .Y(_4031_));
 sky130_fd_sc_hd__a22o_1 _4936_ (.A1(net33),
    .A2(net31),
    .B1(net30),
    .B2(net44),
    .X(_4032_));
 sky130_fd_sc_hd__and4_1 _4937_ (.A(net44),
    .B(net33),
    .C(net30),
    .D(net29),
    .X(_4033_));
 sky130_fd_sc_hd__a22o_1 _4938_ (.A1(net33),
    .A2(net30),
    .B1(net29),
    .B2(net44),
    .X(_4034_));
 sky130_fd_sc_hd__a22oi_2 _4939_ (.A1(net28),
    .A2(net44),
    .B1(net33),
    .B2(net29),
    .Y(_4035_));
 sky130_fd_sc_hd__a22o_1 _4940_ (.A1(net28),
    .A2(net44),
    .B1(net33),
    .B2(net29),
    .X(_4036_));
 sky130_fd_sc_hd__and4_1 _4941_ (.A(net28),
    .B(net44),
    .C(net33),
    .D(net29),
    .X(_4037_));
 sky130_fd_sc_hd__a22oi_2 _4942_ (.A1(net28),
    .A2(net33),
    .B1(net27),
    .B2(net44),
    .Y(_4038_));
 sky130_fd_sc_hd__a22o_1 _4943_ (.A1(net28),
    .A2(net33),
    .B1(net27),
    .B2(net44),
    .X(_4039_));
 sky130_fd_sc_hd__and4_1 _4944_ (.A(net28),
    .B(net44),
    .C(net33),
    .D(net27),
    .X(_4040_));
 sky130_fd_sc_hd__a22o_1 _4945_ (.A1(net33),
    .A2(net27),
    .B1(net26),
    .B2(net44),
    .X(_4041_));
 sky130_fd_sc_hd__and3_1 _4946_ (.A(net44),
    .B(net33),
    .C(net27),
    .X(_4042_));
 sky130_fd_sc_hd__and4_1 _4947_ (.A(net44),
    .B(net33),
    .C(net27),
    .D(net26),
    .X(_4043_));
 sky130_fd_sc_hd__nand2_1 _4948_ (.A(net33),
    .B(net1),
    .Y(_4044_));
 sky130_fd_sc_hd__and4_1 _4949_ (.A(net44),
    .B(net33),
    .C(net12),
    .D(net1),
    .X(_4045_));
 sky130_fd_sc_hd__nand4_1 _4950_ (.A(net44),
    .B(net33),
    .C(net26),
    .D(net23),
    .Y(_4046_));
 sky130_fd_sc_hd__o2111a_1 _4951_ (.A1(net26),
    .A2(net12),
    .B1(net23),
    .C1(net44),
    .D1(net33),
    .X(_4047_));
 sky130_fd_sc_hd__a21o_1 _4952_ (.A1(net26),
    .A2(_4045_),
    .B1(_4047_),
    .X(_4048_));
 sky130_fd_sc_hd__a211o_1 _4953_ (.A1(net26),
    .A2(_4045_),
    .B1(_4047_),
    .C1(_4043_),
    .X(_4049_));
 sky130_fd_sc_hd__a21o_1 _4954_ (.A1(_4041_),
    .A2(_4049_),
    .B1(_4040_),
    .X(_4050_));
 sky130_fd_sc_hd__a21o_1 _4955_ (.A1(_4039_),
    .A2(_4050_),
    .B1(_4037_),
    .X(_4051_));
 sky130_fd_sc_hd__a31o_1 _4956_ (.A1(_4036_),
    .A2(_4039_),
    .A3(_4050_),
    .B1(_4037_),
    .X(_4052_));
 sky130_fd_sc_hd__o211a_2 _4957_ (.A1(_4033_),
    .A2(_4052_),
    .B1(_4034_),
    .C1(_4032_),
    .X(_4053_));
 sky130_fd_sc_hd__o31a_1 _4958_ (.A1(_4028_),
    .A2(_4030_),
    .A3(_4053_),
    .B1(_4029_),
    .X(_4054_));
 sky130_fd_sc_hd__o311ai_4 _4959_ (.A1(_4028_),
    .A2(_4030_),
    .A3(_4053_),
    .B1(_4029_),
    .C1(_4026_),
    .Y(_4055_));
 sky130_fd_sc_hd__a31o_1 _4960_ (.A1(_4025_),
    .A2(_4027_),
    .A3(_4055_),
    .B1(_4023_),
    .X(_4056_));
 sky130_fd_sc_hd__a311o_1 _4961_ (.A1(_4025_),
    .A2(_4027_),
    .A3(_4055_),
    .B1(_4023_),
    .C1(_4022_),
    .X(_4057_));
 sky130_fd_sc_hd__a31o_1 _4962_ (.A1(_4018_),
    .A2(_4020_),
    .A3(_4057_),
    .B1(_4019_),
    .X(_4058_));
 sky130_fd_sc_hd__a311o_1 _4963_ (.A1(_4018_),
    .A2(_4020_),
    .A3(_4057_),
    .B1(_4019_),
    .C1(_4016_),
    .X(_4059_));
 sky130_fd_sc_hd__nand2_1 _4964_ (.A(_4014_),
    .B(_4059_),
    .Y(_4060_));
 sky130_fd_sc_hd__a31oi_2 _4965_ (.A1(_4012_),
    .A2(_4014_),
    .A3(_4059_),
    .B1(_4013_),
    .Y(_4061_));
 sky130_fd_sc_hd__o21a_1 _4966_ (.A1(_4011_),
    .A2(_4061_),
    .B1(_4009_),
    .X(_4062_));
 sky130_fd_sc_hd__o211a_1 _4967_ (.A1(_4011_),
    .A2(_4061_),
    .B1(_4006_),
    .C1(_4009_),
    .X(_4063_));
 sky130_fd_sc_hd__o21bai_1 _4968_ (.A1(_4008_),
    .A2(_4063_),
    .B1_N(_4004_),
    .Y(_4064_));
 sky130_fd_sc_hd__a21o_1 _4969_ (.A1(_4005_),
    .A2(_4064_),
    .B1(_4002_),
    .X(_4065_));
 sky130_fd_sc_hd__a21bo_1 _4970_ (.A1(_4003_),
    .A2(_4065_),
    .B1_N(_4000_),
    .X(_4066_));
 sky130_fd_sc_hd__a31oi_2 _4971_ (.A1(_3998_),
    .A2(_4001_),
    .A3(_4066_),
    .B1(_3999_),
    .Y(_4067_));
 sky130_fd_sc_hd__o21ai_1 _4972_ (.A1(_3995_),
    .A2(_4067_),
    .B1(_3996_),
    .Y(_4068_));
 sky130_fd_sc_hd__o211a_1 _4973_ (.A1(_3995_),
    .A2(_4067_),
    .B1(_3996_),
    .C1(_3994_),
    .X(_4069_));
 sky130_fd_sc_hd__a21oi_2 _4974_ (.A1(_1716_),
    .A2(_4069_),
    .B1(_3993_),
    .Y(_4070_));
 sky130_fd_sc_hd__a21o_1 _4975_ (.A1(net44),
    .A2(_1716_),
    .B1(_4069_),
    .X(_4071_));
 sky130_fd_sc_hd__a22o_1 _4976_ (.A1(net55),
    .A2(net15),
    .B1(_4070_),
    .B2(_4071_),
    .X(_4072_));
 sky130_fd_sc_hd__and4_1 _4977_ (.A(net55),
    .B(net15),
    .C(_4070_),
    .D(_4071_),
    .X(_4073_));
 sky130_fd_sc_hd__nand4_1 _4978_ (.A(net55),
    .B(net15),
    .C(_4070_),
    .D(_4071_),
    .Y(_4074_));
 sky130_fd_sc_hd__and2_1 _4979_ (.A(net55),
    .B(net14),
    .X(_4075_));
 sky130_fd_sc_hd__and2b_1 _4980_ (.A_N(_3993_),
    .B(_3994_),
    .X(_4076_));
 sky130_fd_sc_hd__xnor2_1 _4981_ (.A(_4068_),
    .B(_4076_),
    .Y(_4077_));
 sky130_fd_sc_hd__and2_1 _4982_ (.A(_4075_),
    .B(_4077_),
    .X(_4078_));
 sky130_fd_sc_hd__nand2_1 _4983_ (.A(net55),
    .B(net13),
    .Y(_4079_));
 sky130_fd_sc_hd__nand2b_1 _4984_ (.A_N(_3995_),
    .B(_3996_),
    .Y(_4080_));
 sky130_fd_sc_hd__xnor2_1 _4985_ (.A(_4067_),
    .B(_4080_),
    .Y(_4081_));
 sky130_fd_sc_hd__and3_1 _4986_ (.A(net55),
    .B(net13),
    .C(_4081_),
    .X(_4082_));
 sky130_fd_sc_hd__a21o_1 _4987_ (.A1(net55),
    .A2(net13),
    .B1(_4081_),
    .X(_4083_));
 sky130_fd_sc_hd__nand2_1 _4988_ (.A(net55),
    .B(net11),
    .Y(_4084_));
 sky130_fd_sc_hd__nor2_1 _4989_ (.A(_3997_),
    .B(_3999_),
    .Y(_4085_));
 sky130_fd_sc_hd__a21o_1 _4990_ (.A1(_4001_),
    .A2(_4066_),
    .B1(_4085_),
    .X(_4086_));
 sky130_fd_sc_hd__nand3_1 _4991_ (.A(_4001_),
    .B(_4066_),
    .C(_4085_),
    .Y(_4087_));
 sky130_fd_sc_hd__and3_1 _4992_ (.A(_4084_),
    .B(_4086_),
    .C(_4087_),
    .X(_4088_));
 sky130_fd_sc_hd__nand3_1 _4993_ (.A(_4084_),
    .B(_4086_),
    .C(_4087_),
    .Y(_4089_));
 sky130_fd_sc_hd__a21oi_1 _4994_ (.A1(_4086_),
    .A2(_4087_),
    .B1(_4084_),
    .Y(_4090_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_4000_),
    .B(_4001_),
    .Y(_4091_));
 sky130_fd_sc_hd__nand3_1 _4996_ (.A(_4003_),
    .B(_4065_),
    .C(_4091_),
    .Y(_4092_));
 sky130_fd_sc_hd__a21o_1 _4997_ (.A1(_4003_),
    .A2(_4065_),
    .B1(_4091_),
    .X(_4093_));
 sky130_fd_sc_hd__and4_1 _4998_ (.A(net55),
    .B(net10),
    .C(_4092_),
    .D(_4093_),
    .X(_4094_));
 sky130_fd_sc_hd__a22oi_2 _4999_ (.A1(net55),
    .A2(net10),
    .B1(_4092_),
    .B2(_4093_),
    .Y(_4095_));
 sky130_fd_sc_hd__nand2b_1 _5000_ (.A_N(_4002_),
    .B(_4003_),
    .Y(_4096_));
 sky130_fd_sc_hd__nand3_1 _5001_ (.A(_4005_),
    .B(_4064_),
    .C(_4096_),
    .Y(_4097_));
 sky130_fd_sc_hd__a21o_1 _5002_ (.A1(_4005_),
    .A2(_4064_),
    .B1(_4096_),
    .X(_4098_));
 sky130_fd_sc_hd__and4_1 _5003_ (.A(net55),
    .B(net9),
    .C(_4097_),
    .D(_4098_),
    .X(_4099_));
 sky130_fd_sc_hd__nand4_1 _5004_ (.A(net55),
    .B(net9),
    .C(_4097_),
    .D(_4098_),
    .Y(_4100_));
 sky130_fd_sc_hd__a22o_1 _5005_ (.A1(net55),
    .A2(net9),
    .B1(_4097_),
    .B2(_4098_),
    .X(_4101_));
 sky130_fd_sc_hd__and2_1 _5006_ (.A(net55),
    .B(net8),
    .X(_4102_));
 sky130_fd_sc_hd__and2b_1 _5007_ (.A_N(_4004_),
    .B(_4005_),
    .X(_4103_));
 sky130_fd_sc_hd__or3_1 _5008_ (.A(_4008_),
    .B(_4063_),
    .C(_4103_),
    .X(_4104_));
 sky130_fd_sc_hd__o21ai_1 _5009_ (.A1(_4008_),
    .A2(_4063_),
    .B1(_4103_),
    .Y(_4105_));
 sky130_fd_sc_hd__and2_1 _5010_ (.A(_4104_),
    .B(_4105_),
    .X(_4106_));
 sky130_fd_sc_hd__a21o_1 _5011_ (.A1(_4104_),
    .A2(_4105_),
    .B1(_4102_),
    .X(_4107_));
 sky130_fd_sc_hd__and3_1 _5012_ (.A(_4102_),
    .B(_4104_),
    .C(_4105_),
    .X(_4108_));
 sky130_fd_sc_hd__nand2_1 _5013_ (.A(net55),
    .B(net7),
    .Y(_4109_));
 sky130_fd_sc_hd__a21bo_1 _5014_ (.A1(net9),
    .A2(_4007_),
    .B1_N(_4006_),
    .X(_4110_));
 sky130_fd_sc_hd__xnor2_1 _5015_ (.A(_4062_),
    .B(_4110_),
    .Y(_4111_));
 sky130_fd_sc_hd__nand2b_1 _5016_ (.A_N(_4111_),
    .B(_4109_),
    .Y(_4112_));
 sky130_fd_sc_hd__and3_1 _5017_ (.A(net55),
    .B(net7),
    .C(_4111_),
    .X(_4113_));
 sky130_fd_sc_hd__nand2_1 _5018_ (.A(net55),
    .B(net6),
    .Y(_4114_));
 sky130_fd_sc_hd__a21boi_1 _5019_ (.A1(net8),
    .A2(_4010_),
    .B1_N(_4009_),
    .Y(_4115_));
 sky130_fd_sc_hd__xnor2_1 _5020_ (.A(_4061_),
    .B(_4115_),
    .Y(_4116_));
 sky130_fd_sc_hd__and2_1 _5021_ (.A(_4114_),
    .B(_4116_),
    .X(_4117_));
 sky130_fd_sc_hd__nor2_1 _5022_ (.A(_4114_),
    .B(_4116_),
    .Y(_4118_));
 sky130_fd_sc_hd__nand2_1 _5023_ (.A(net55),
    .B(net5),
    .Y(_4119_));
 sky130_fd_sc_hd__a21o_1 _5024_ (.A1(net6),
    .A2(_4010_),
    .B1(_4013_),
    .X(_4120_));
 sky130_fd_sc_hd__xnor2_1 _5025_ (.A(_4060_),
    .B(_4120_),
    .Y(_4121_));
 sky130_fd_sc_hd__nand2b_1 _5026_ (.A_N(_4119_),
    .B(_4121_),
    .Y(_4122_));
 sky130_fd_sc_hd__a21oi_1 _5027_ (.A1(net55),
    .A2(net5),
    .B1(_4121_),
    .Y(_4123_));
 sky130_fd_sc_hd__nand2_1 _5028_ (.A(net55),
    .B(net4),
    .Y(_4124_));
 sky130_fd_sc_hd__nand2_1 _5029_ (.A(_4014_),
    .B(_4015_),
    .Y(_4125_));
 sky130_fd_sc_hd__xor2_1 _5030_ (.A(_4058_),
    .B(_4125_),
    .X(_4126_));
 sky130_fd_sc_hd__nand2b_1 _5031_ (.A_N(_4124_),
    .B(_4126_),
    .Y(_4127_));
 sky130_fd_sc_hd__a21oi_1 _5032_ (.A1(net55),
    .A2(net4),
    .B1(_4126_),
    .Y(_4128_));
 sky130_fd_sc_hd__nand2_1 _5033_ (.A(net55),
    .B(net3),
    .Y(_4129_));
 sky130_fd_sc_hd__nor2_1 _5034_ (.A(_4017_),
    .B(_4019_),
    .Y(_4130_));
 sky130_fd_sc_hd__a21o_1 _5035_ (.A1(_4020_),
    .A2(_4057_),
    .B1(_4130_),
    .X(_4131_));
 sky130_fd_sc_hd__nand3_1 _5036_ (.A(_4020_),
    .B(_4057_),
    .C(_4130_),
    .Y(_4132_));
 sky130_fd_sc_hd__and3_1 _5037_ (.A(_4129_),
    .B(_4131_),
    .C(_4132_),
    .X(_4133_));
 sky130_fd_sc_hd__a21o_1 _5038_ (.A1(_4131_),
    .A2(_4132_),
    .B1(_4129_),
    .X(_4134_));
 sky130_fd_sc_hd__nand2_1 _5039_ (.A(net55),
    .B(net2),
    .Y(_4135_));
 sky130_fd_sc_hd__nand2_1 _5040_ (.A(_4020_),
    .B(_4021_),
    .Y(_4136_));
 sky130_fd_sc_hd__xor2_1 _5041_ (.A(_4056_),
    .B(_4136_),
    .X(_4137_));
 sky130_fd_sc_hd__a21oi_1 _5042_ (.A1(net55),
    .A2(net2),
    .B1(_4137_),
    .Y(_4138_));
 sky130_fd_sc_hd__nand2b_1 _5043_ (.A_N(_4135_),
    .B(_4137_),
    .Y(_4139_));
 sky130_fd_sc_hd__nand2_1 _5044_ (.A(net55),
    .B(net32),
    .Y(_4140_));
 sky130_fd_sc_hd__nor2_1 _5045_ (.A(_4023_),
    .B(_4024_),
    .Y(_4141_));
 sky130_fd_sc_hd__a21o_1 _5046_ (.A1(_4027_),
    .A2(_4055_),
    .B1(_4141_),
    .X(_4142_));
 sky130_fd_sc_hd__nand3_1 _5047_ (.A(_4027_),
    .B(_4055_),
    .C(_4141_),
    .Y(_4143_));
 sky130_fd_sc_hd__a21oi_2 _5048_ (.A1(_4142_),
    .A2(_4143_),
    .B1(_4140_),
    .Y(_4144_));
 sky130_fd_sc_hd__inv_2 _5049_ (.A(_4144_),
    .Y(_4145_));
 sky130_fd_sc_hd__and3_1 _5050_ (.A(_4140_),
    .B(_4142_),
    .C(_4143_),
    .X(_4146_));
 sky130_fd_sc_hd__nand3_1 _5051_ (.A(_4140_),
    .B(_4142_),
    .C(_4143_),
    .Y(_4147_));
 sky130_fd_sc_hd__nand2_2 _5052_ (.A(net55),
    .B(net31),
    .Y(_4148_));
 sky130_fd_sc_hd__nand2_1 _5053_ (.A(_4026_),
    .B(_4027_),
    .Y(_4149_));
 sky130_fd_sc_hd__xor2_2 _5054_ (.A(_4054_),
    .B(_4149_),
    .X(_4150_));
 sky130_fd_sc_hd__nand2_1 _5055_ (.A(_4148_),
    .B(_4150_),
    .Y(_4151_));
 sky130_fd_sc_hd__nand2_1 _5056_ (.A(net55),
    .B(net30),
    .Y(_4152_));
 sky130_fd_sc_hd__and2b_1 _5057_ (.A_N(_4028_),
    .B(_4029_),
    .X(_4153_));
 sky130_fd_sc_hd__o21bai_1 _5058_ (.A1(_4030_),
    .A2(_4053_),
    .B1_N(_4153_),
    .Y(_4154_));
 sky130_fd_sc_hd__or3b_1 _5059_ (.A(_4030_),
    .B(_4053_),
    .C_N(_4153_),
    .X(_4155_));
 sky130_fd_sc_hd__and3_1 _5060_ (.A(_4152_),
    .B(_4154_),
    .C(_4155_),
    .X(_4156_));
 sky130_fd_sc_hd__nand3_1 _5061_ (.A(_4152_),
    .B(_4154_),
    .C(_4155_),
    .Y(_4157_));
 sky130_fd_sc_hd__a21o_1 _5062_ (.A1(_4154_),
    .A2(_4155_),
    .B1(_4152_),
    .X(_4158_));
 sky130_fd_sc_hd__and2_1 _5063_ (.A(_4031_),
    .B(_4032_),
    .X(_4159_));
 sky130_fd_sc_hd__a311o_1 _5064_ (.A1(_4034_),
    .A2(_4036_),
    .A3(_4051_),
    .B1(_4159_),
    .C1(_4033_),
    .X(_4160_));
 sky130_fd_sc_hd__o211ai_2 _5065_ (.A1(_4033_),
    .A2(_4052_),
    .B1(_4159_),
    .C1(_4034_),
    .Y(_4161_));
 sky130_fd_sc_hd__a22oi_2 _5066_ (.A1(net55),
    .A2(net29),
    .B1(_4160_),
    .B2(_4161_),
    .Y(_4162_));
 sky130_fd_sc_hd__a22o_1 _5067_ (.A1(net55),
    .A2(net29),
    .B1(_4160_),
    .B2(_4161_),
    .X(_4163_));
 sky130_fd_sc_hd__and4_1 _5068_ (.A(net55),
    .B(net29),
    .C(_4160_),
    .D(_4161_),
    .X(_4164_));
 sky130_fd_sc_hd__nand2_1 _5069_ (.A(net28),
    .B(net55),
    .Y(_4165_));
 sky130_fd_sc_hd__inv_2 _5070_ (.A(_4165_),
    .Y(_4166_));
 sky130_fd_sc_hd__nand2b_1 _5071_ (.A_N(_4033_),
    .B(_4034_),
    .Y(_4167_));
 sky130_fd_sc_hd__xnor2_1 _5072_ (.A(_4052_),
    .B(_4167_),
    .Y(_4168_));
 sky130_fd_sc_hd__and2_1 _5073_ (.A(_4166_),
    .B(_4168_),
    .X(_4169_));
 sky130_fd_sc_hd__nand2_1 _5074_ (.A(net27),
    .B(net55),
    .Y(_4170_));
 sky130_fd_sc_hd__a211o_1 _5075_ (.A1(_4039_),
    .A2(_4050_),
    .B1(_4035_),
    .C1(_4037_),
    .X(_4171_));
 sky130_fd_sc_hd__o211ai_2 _5076_ (.A1(_4035_),
    .A2(_4037_),
    .B1(_4039_),
    .C1(_4050_),
    .Y(_4172_));
 sky130_fd_sc_hd__a21oi_1 _5077_ (.A1(_4171_),
    .A2(_4172_),
    .B1(_4170_),
    .Y(_4173_));
 sky130_fd_sc_hd__a21o_1 _5078_ (.A1(_4171_),
    .A2(_4172_),
    .B1(_4170_),
    .X(_4174_));
 sky130_fd_sc_hd__and3_1 _5079_ (.A(_4170_),
    .B(_4171_),
    .C(_4172_),
    .X(_4175_));
 sky130_fd_sc_hd__nand3_1 _5080_ (.A(_4170_),
    .B(_4171_),
    .C(_4172_),
    .Y(_4176_));
 sky130_fd_sc_hd__nand2_1 _5081_ (.A(net26),
    .B(net55),
    .Y(_4177_));
 sky130_fd_sc_hd__o211ai_2 _5082_ (.A1(_4038_),
    .A2(_4040_),
    .B1(_4041_),
    .C1(_4049_),
    .Y(_4178_));
 sky130_fd_sc_hd__a211o_1 _5083_ (.A1(_4041_),
    .A2(_4049_),
    .B1(_4038_),
    .C1(_4040_),
    .X(_4179_));
 sky130_fd_sc_hd__and3_1 _5084_ (.A(_4177_),
    .B(_4178_),
    .C(_4179_),
    .X(_4180_));
 sky130_fd_sc_hd__nand3_1 _5085_ (.A(_4177_),
    .B(_4178_),
    .C(_4179_),
    .Y(_4181_));
 sky130_fd_sc_hd__a21oi_1 _5086_ (.A1(_4178_),
    .A2(_4179_),
    .B1(_4177_),
    .Y(_4182_));
 sky130_fd_sc_hd__nand2_1 _5087_ (.A(net23),
    .B(net55),
    .Y(_4183_));
 sky130_fd_sc_hd__inv_2 _5088_ (.A(_4183_),
    .Y(_4184_));
 sky130_fd_sc_hd__a21bo_1 _5089_ (.A1(net26),
    .A2(_4042_),
    .B1_N(_4041_),
    .X(_4185_));
 sky130_fd_sc_hd__xnor2_1 _5090_ (.A(_4048_),
    .B(_4185_),
    .Y(_4186_));
 sky130_fd_sc_hd__or2_1 _5091_ (.A(_4184_),
    .B(_4186_),
    .X(_4188_));
 sky130_fd_sc_hd__a22o_1 _5092_ (.A1(net33),
    .A2(net26),
    .B1(net23),
    .B2(net44),
    .X(_4189_));
 sky130_fd_sc_hd__o2111a_1 _5093_ (.A1(net23),
    .A2(net1),
    .B1(net12),
    .C1(net44),
    .D1(net33),
    .X(_4190_));
 sky130_fd_sc_hd__nand3_1 _5094_ (.A(_4046_),
    .B(_4189_),
    .C(_4190_),
    .Y(_4191_));
 sky130_fd_sc_hd__a21o_1 _5095_ (.A1(_4046_),
    .A2(_4189_),
    .B1(_4190_),
    .X(_4192_));
 sky130_fd_sc_hd__and4_1 _5096_ (.A(net12),
    .B(net55),
    .C(_4191_),
    .D(_4192_),
    .X(_4193_));
 sky130_fd_sc_hd__nand4_1 _5097_ (.A(net12),
    .B(net55),
    .C(_4191_),
    .D(_4192_),
    .Y(_4194_));
 sky130_fd_sc_hd__a22o_1 _5098_ (.A1(net12),
    .A2(net55),
    .B1(_4191_),
    .B2(_4192_),
    .X(_4195_));
 sky130_fd_sc_hd__a32o_1 _5099_ (.A1(net44),
    .A2(net12),
    .A3(_4044_),
    .B1(net33),
    .B2(net23),
    .X(_4196_));
 sky130_fd_sc_hd__and3_1 _5100_ (.A(net1),
    .B(net55),
    .C(_4196_),
    .X(_4197_));
 sky130_fd_sc_hd__a21oi_1 _5101_ (.A1(_4195_),
    .A2(_4197_),
    .B1(_4193_),
    .Y(_4199_));
 sky130_fd_sc_hd__a221o_1 _5102_ (.A1(_4184_),
    .A2(_4186_),
    .B1(_4195_),
    .B2(_4197_),
    .C1(_4193_),
    .X(_4200_));
 sky130_fd_sc_hd__a31o_1 _5103_ (.A1(_4181_),
    .A2(_4188_),
    .A3(_4200_),
    .B1(_4182_),
    .X(_4201_));
 sky130_fd_sc_hd__a31oi_1 _5104_ (.A1(_4181_),
    .A2(_4188_),
    .A3(_4200_),
    .B1(_4182_),
    .Y(_4202_));
 sky130_fd_sc_hd__a21oi_1 _5105_ (.A1(_4174_),
    .A2(_4202_),
    .B1(_4175_),
    .Y(_4203_));
 sky130_fd_sc_hd__o221a_2 _5106_ (.A1(_4166_),
    .A2(_4168_),
    .B1(_4173_),
    .B2(_4201_),
    .C1(_4176_),
    .X(_4204_));
 sky130_fd_sc_hd__o31ai_4 _5107_ (.A1(_4164_),
    .A2(_4169_),
    .A3(_4204_),
    .B1(_4163_),
    .Y(_4205_));
 sky130_fd_sc_hd__o21a_1 _5108_ (.A1(_4156_),
    .A2(_4205_),
    .B1(_4158_),
    .X(_4206_));
 sky130_fd_sc_hd__o221ai_4 _5109_ (.A1(_4148_),
    .A2(_4150_),
    .B1(_4156_),
    .B2(_4205_),
    .C1(_4158_),
    .Y(_4207_));
 sky130_fd_sc_hd__nand3_1 _5110_ (.A(_4147_),
    .B(_4151_),
    .C(_4207_),
    .Y(_4208_));
 sky130_fd_sc_hd__a21o_1 _5111_ (.A1(_4151_),
    .A2(_4207_),
    .B1(_4144_),
    .X(_0001_));
 sky130_fd_sc_hd__a31o_1 _5112_ (.A1(_4139_),
    .A2(_4145_),
    .A3(_4208_),
    .B1(_4138_),
    .X(_0002_));
 sky130_fd_sc_hd__a311o_1 _5113_ (.A1(_4139_),
    .A2(_4145_),
    .A3(_4208_),
    .B1(_4138_),
    .C1(_4133_),
    .X(_0003_));
 sky130_fd_sc_hd__a31o_1 _5114_ (.A1(_4127_),
    .A2(_4134_),
    .A3(_0003_),
    .B1(_4128_),
    .X(_0004_));
 sky130_fd_sc_hd__a21oi_1 _5115_ (.A1(_4122_),
    .A2(_0004_),
    .B1(_4123_),
    .Y(_0005_));
 sky130_fd_sc_hd__a211oi_2 _5116_ (.A1(_4122_),
    .A2(_0004_),
    .B1(_4123_),
    .C1(_4117_),
    .Y(_0006_));
 sky130_fd_sc_hd__o31a_1 _5117_ (.A1(_4113_),
    .A2(_4118_),
    .A3(_0006_),
    .B1(_4112_),
    .X(_0007_));
 sky130_fd_sc_hd__o311a_1 _5118_ (.A1(_4113_),
    .A2(_4118_),
    .A3(_0006_),
    .B1(_4112_),
    .C1(_4107_),
    .X(_0008_));
 sky130_fd_sc_hd__o31ai_1 _5119_ (.A1(_4099_),
    .A2(_4108_),
    .A3(_0008_),
    .B1(_4101_),
    .Y(_0009_));
 sky130_fd_sc_hd__o31a_1 _5120_ (.A1(_4099_),
    .A2(_4108_),
    .A3(_0008_),
    .B1(_4101_),
    .X(_0010_));
 sky130_fd_sc_hd__o21ba_1 _5121_ (.A1(_4094_),
    .A2(_0010_),
    .B1_N(_4095_),
    .X(_0012_));
 sky130_fd_sc_hd__a21o_1 _5122_ (.A1(_4089_),
    .A2(_0012_),
    .B1(_4090_),
    .X(_0013_));
 sky130_fd_sc_hd__o21ai_1 _5123_ (.A1(_4082_),
    .A2(_0013_),
    .B1(_4083_),
    .Y(_0014_));
 sky130_fd_sc_hd__o221a_1 _5124_ (.A1(_4075_),
    .A2(_4077_),
    .B1(_4082_),
    .B2(_0013_),
    .C1(_4083_),
    .X(_0015_));
 sky130_fd_sc_hd__o31a_1 _5125_ (.A1(_4073_),
    .A2(_4078_),
    .A3(_0015_),
    .B1(_4072_),
    .X(_0016_));
 sky130_fd_sc_hd__o311a_1 _5126_ (.A1(_3993_),
    .A2(_4069_),
    .A3(_0016_),
    .B1(_1716_),
    .C1(net55),
    .X(_0017_));
 sky130_fd_sc_hd__nor2_1 _5127_ (.A(_0022_),
    .B(_1727_),
    .Y(_0018_));
 sky130_fd_sc_hd__mux2_1 _5128_ (.A0(_0018_),
    .A1(_0022_),
    .S(_0017_),
    .X(_0019_));
 sky130_fd_sc_hd__xnor2_1 _5129_ (.A(_4070_),
    .B(_0016_),
    .Y(_0020_));
 sky130_fd_sc_hd__xnor2_1 _5130_ (.A(_3991_),
    .B(_0020_),
    .Y(_0021_));
 sky130_fd_sc_hd__a211o_1 _5131_ (.A1(_4072_),
    .A2(_4074_),
    .B1(_4078_),
    .C1(_0015_),
    .X(_0023_));
 sky130_fd_sc_hd__o211ai_2 _5132_ (.A1(_4078_),
    .A2(_0015_),
    .B1(_4072_),
    .C1(_4074_),
    .Y(_0024_));
 sky130_fd_sc_hd__a22o_1 _5133_ (.A1(net14),
    .A2(net58),
    .B1(_0023_),
    .B2(_0024_),
    .X(_0025_));
 sky130_fd_sc_hd__and4_1 _5134_ (.A(net14),
    .B(net58),
    .C(_0023_),
    .D(_0024_),
    .X(_0026_));
 sky130_fd_sc_hd__nand4_1 _5135_ (.A(net14),
    .B(net58),
    .C(_0023_),
    .D(_0024_),
    .Y(_0027_));
 sky130_fd_sc_hd__nand2_1 _5136_ (.A(net13),
    .B(net58),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _5137_ (.A(_0028_),
    .Y(_0029_));
 sky130_fd_sc_hd__xor2_1 _5138_ (.A(_4075_),
    .B(_4077_),
    .X(_0030_));
 sky130_fd_sc_hd__xnor2_1 _5139_ (.A(_0014_),
    .B(_0030_),
    .Y(_0031_));
 sky130_fd_sc_hd__and2_1 _5140_ (.A(_0029_),
    .B(_0031_),
    .X(_0032_));
 sky130_fd_sc_hd__xor2_1 _5141_ (.A(_4079_),
    .B(_4081_),
    .X(_0034_));
 sky130_fd_sc_hd__xnor2_1 _5142_ (.A(_0013_),
    .B(_0034_),
    .Y(_0035_));
 sky130_fd_sc_hd__and2_1 _5143_ (.A(net11),
    .B(net58),
    .X(_0036_));
 sky130_fd_sc_hd__or2_1 _5144_ (.A(_0035_),
    .B(_0036_),
    .X(_0037_));
 sky130_fd_sc_hd__nand2_1 _5145_ (.A(net10),
    .B(net58),
    .Y(_0038_));
 sky130_fd_sc_hd__o21ai_1 _5146_ (.A1(_4088_),
    .A2(_4090_),
    .B1(_0012_),
    .Y(_0039_));
 sky130_fd_sc_hd__or3_1 _5147_ (.A(_4088_),
    .B(_4090_),
    .C(_0012_),
    .X(_0040_));
 sky130_fd_sc_hd__nand3_1 _5148_ (.A(_0038_),
    .B(_0039_),
    .C(_0040_),
    .Y(_0041_));
 sky130_fd_sc_hd__a21oi_1 _5149_ (.A1(_0039_),
    .A2(_0040_),
    .B1(_0038_),
    .Y(_0042_));
 sky130_fd_sc_hd__a21o_1 _5150_ (.A1(_0039_),
    .A2(_0040_),
    .B1(_0038_),
    .X(_0043_));
 sky130_fd_sc_hd__o21ai_1 _5151_ (.A1(_4094_),
    .A2(_4095_),
    .B1(_0009_),
    .Y(_0045_));
 sky130_fd_sc_hd__or3_1 _5152_ (.A(_4094_),
    .B(_4095_),
    .C(_0009_),
    .X(_0046_));
 sky130_fd_sc_hd__and4_1 _5153_ (.A(net9),
    .B(net58),
    .C(_0045_),
    .D(_0046_),
    .X(_0047_));
 sky130_fd_sc_hd__a22oi_2 _5154_ (.A1(net9),
    .A2(net58),
    .B1(_0045_),
    .B2(_0046_),
    .Y(_0048_));
 sky130_fd_sc_hd__a22o_1 _5155_ (.A1(net9),
    .A2(net58),
    .B1(_0045_),
    .B2(_0046_),
    .X(_0049_));
 sky130_fd_sc_hd__and2_1 _5156_ (.A(net8),
    .B(net58),
    .X(_0050_));
 sky130_fd_sc_hd__a211o_1 _5157_ (.A1(_4100_),
    .A2(_4101_),
    .B1(_4108_),
    .C1(_0008_),
    .X(_0051_));
 sky130_fd_sc_hd__o211ai_2 _5158_ (.A1(_4108_),
    .A2(_0008_),
    .B1(_4100_),
    .C1(_4101_),
    .Y(_0052_));
 sky130_fd_sc_hd__a21oi_1 _5159_ (.A1(_0051_),
    .A2(_0052_),
    .B1(_0050_),
    .Y(_0053_));
 sky130_fd_sc_hd__a21o_1 _5160_ (.A1(_0051_),
    .A2(_0052_),
    .B1(_0050_),
    .X(_0054_));
 sky130_fd_sc_hd__and3_1 _5161_ (.A(_0050_),
    .B(_0051_),
    .C(_0052_),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_1 _5162_ (.A(net7),
    .B(net58),
    .Y(_0057_));
 sky130_fd_sc_hd__xor2_1 _5163_ (.A(_4102_),
    .B(_4106_),
    .X(_0058_));
 sky130_fd_sc_hd__xor2_1 _5164_ (.A(_0007_),
    .B(_0058_),
    .X(_0059_));
 sky130_fd_sc_hd__a21o_1 _5165_ (.A1(net7),
    .A2(net58),
    .B1(_0059_),
    .X(_0060_));
 sky130_fd_sc_hd__and3_1 _5166_ (.A(net7),
    .B(net58),
    .C(_0059_),
    .X(_0061_));
 sky130_fd_sc_hd__xor2_1 _5167_ (.A(_4109_),
    .B(_4111_),
    .X(_0062_));
 sky130_fd_sc_hd__or3b_1 _5168_ (.A(_4118_),
    .B(_0006_),
    .C_N(_0062_),
    .X(_0063_));
 sky130_fd_sc_hd__o21bai_1 _5169_ (.A1(_4118_),
    .A2(_0006_),
    .B1_N(_0062_),
    .Y(_0064_));
 sky130_fd_sc_hd__and4_1 _5170_ (.A(net6),
    .B(net58),
    .C(_0063_),
    .D(_0064_),
    .X(_0065_));
 sky130_fd_sc_hd__a22o_1 _5171_ (.A1(net6),
    .A2(net58),
    .B1(_0063_),
    .B2(_0064_),
    .X(_0067_));
 sky130_fd_sc_hd__nand2_1 _5172_ (.A(net5),
    .B(net58),
    .Y(_0068_));
 sky130_fd_sc_hd__nor2_1 _5173_ (.A(_4117_),
    .B(_4118_),
    .Y(_0069_));
 sky130_fd_sc_hd__xnor2_1 _5174_ (.A(_0005_),
    .B(_0069_),
    .Y(_0070_));
 sky130_fd_sc_hd__nand2_1 _5175_ (.A(_0068_),
    .B(_0070_),
    .Y(_0071_));
 sky130_fd_sc_hd__nor2_1 _5176_ (.A(_0068_),
    .B(_0070_),
    .Y(_0072_));
 sky130_fd_sc_hd__nand2_1 _5177_ (.A(net4),
    .B(net58),
    .Y(_0073_));
 sky130_fd_sc_hd__xnor2_1 _5178_ (.A(_4119_),
    .B(_4121_),
    .Y(_0074_));
 sky130_fd_sc_hd__xnor2_1 _5179_ (.A(_0004_),
    .B(_0074_),
    .Y(_0075_));
 sky130_fd_sc_hd__nand2b_1 _5180_ (.A_N(_0075_),
    .B(_0073_),
    .Y(_0076_));
 sky130_fd_sc_hd__and3_1 _5181_ (.A(net4),
    .B(net58),
    .C(_0075_),
    .X(_0078_));
 sky130_fd_sc_hd__nand2_1 _5182_ (.A(net3),
    .B(net58),
    .Y(_0079_));
 sky130_fd_sc_hd__xnor2_1 _5183_ (.A(_4124_),
    .B(_4126_),
    .Y(_0080_));
 sky130_fd_sc_hd__nand3_1 _5184_ (.A(_4134_),
    .B(_0003_),
    .C(_0080_),
    .Y(_0081_));
 sky130_fd_sc_hd__a21o_1 _5185_ (.A1(_4134_),
    .A2(_0003_),
    .B1(_0080_),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _5186_ (.A(_0081_),
    .B(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__a21o_1 _5187_ (.A1(_0081_),
    .A2(_0082_),
    .B1(_0079_),
    .X(_0084_));
 sky130_fd_sc_hd__nand2_1 _5188_ (.A(_0079_),
    .B(_0083_),
    .Y(_0085_));
 sky130_fd_sc_hd__nand2_1 _5189_ (.A(net2),
    .B(net58),
    .Y(_0086_));
 sky130_fd_sc_hd__and2b_1 _5190_ (.A_N(_4133_),
    .B(_4134_),
    .X(_0087_));
 sky130_fd_sc_hd__xnor2_1 _5191_ (.A(_0002_),
    .B(_0087_),
    .Y(_0089_));
 sky130_fd_sc_hd__a21oi_1 _5192_ (.A1(net2),
    .A2(net58),
    .B1(_0089_),
    .Y(_0090_));
 sky130_fd_sc_hd__nand2b_1 _5193_ (.A_N(_0086_),
    .B(_0089_),
    .Y(_0091_));
 sky130_fd_sc_hd__nand2_1 _5194_ (.A(net32),
    .B(net58),
    .Y(_0092_));
 sky130_fd_sc_hd__xor2_1 _5195_ (.A(_4135_),
    .B(_4137_),
    .X(_0093_));
 sky130_fd_sc_hd__nand3_1 _5196_ (.A(_4147_),
    .B(_0001_),
    .C(_0093_),
    .Y(_0094_));
 sky130_fd_sc_hd__a21o_1 _5197_ (.A1(_4147_),
    .A2(_0001_),
    .B1(_0093_),
    .X(_0095_));
 sky130_fd_sc_hd__nand3_1 _5198_ (.A(_0092_),
    .B(_0094_),
    .C(_0095_),
    .Y(_0096_));
 sky130_fd_sc_hd__a21o_1 _5199_ (.A1(_0094_),
    .A2(_0095_),
    .B1(_0092_),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _5200_ (.A(net31),
    .B(net58),
    .X(_0098_));
 sky130_fd_sc_hd__a2bb2o_1 _5201_ (.A1_N(_4144_),
    .A2_N(_4146_),
    .B1(_4151_),
    .B2(_4207_),
    .X(_0100_));
 sky130_fd_sc_hd__or4bb_1 _5202_ (.A(_4144_),
    .B(_4146_),
    .C_N(_4151_),
    .D_N(_4207_),
    .X(_0101_));
 sky130_fd_sc_hd__a21oi_1 _5203_ (.A1(_0100_),
    .A2(_0101_),
    .B1(_0098_),
    .Y(_0102_));
 sky130_fd_sc_hd__a21o_1 _5204_ (.A1(_0100_),
    .A2(_0101_),
    .B1(_0098_),
    .X(_0103_));
 sky130_fd_sc_hd__and3_1 _5205_ (.A(_0098_),
    .B(_0100_),
    .C(_0101_),
    .X(_0104_));
 sky130_fd_sc_hd__nand2_1 _5206_ (.A(net30),
    .B(net58),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _5207_ (.A(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hd__xor2_1 _5208_ (.A(_4148_),
    .B(_4150_),
    .X(_0107_));
 sky130_fd_sc_hd__xnor2_1 _5209_ (.A(_4206_),
    .B(_0107_),
    .Y(_0108_));
 sky130_fd_sc_hd__and2_1 _5210_ (.A(_0106_),
    .B(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__nand2_1 _5211_ (.A(net29),
    .B(net58),
    .Y(_0111_));
 sky130_fd_sc_hd__a21o_1 _5212_ (.A1(_4157_),
    .A2(_4158_),
    .B1(_4205_),
    .X(_0112_));
 sky130_fd_sc_hd__nand3_1 _5213_ (.A(_4157_),
    .B(_4158_),
    .C(_4205_),
    .Y(_0113_));
 sky130_fd_sc_hd__a21oi_1 _5214_ (.A1(_0112_),
    .A2(_0113_),
    .B1(_0111_),
    .Y(_0114_));
 sky130_fd_sc_hd__a21o_1 _5215_ (.A1(_0112_),
    .A2(_0113_),
    .B1(_0111_),
    .X(_0115_));
 sky130_fd_sc_hd__and3_1 _5216_ (.A(_0111_),
    .B(_0112_),
    .C(_0113_),
    .X(_0116_));
 sky130_fd_sc_hd__nand3_1 _5217_ (.A(_0111_),
    .B(_0112_),
    .C(_0113_),
    .Y(_0117_));
 sky130_fd_sc_hd__nand2_1 _5218_ (.A(net28),
    .B(net58),
    .Y(_0118_));
 sky130_fd_sc_hd__o22ai_2 _5219_ (.A1(_4162_),
    .A2(_4164_),
    .B1(_4169_),
    .B2(_4204_),
    .Y(_0119_));
 sky130_fd_sc_hd__or4_1 _5220_ (.A(_4162_),
    .B(_4164_),
    .C(_4169_),
    .D(_4204_),
    .X(_0120_));
 sky130_fd_sc_hd__a21oi_1 _5221_ (.A1(_0119_),
    .A2(_0120_),
    .B1(_0118_),
    .Y(_0122_));
 sky130_fd_sc_hd__a21o_1 _5222_ (.A1(_0119_),
    .A2(_0120_),
    .B1(_0118_),
    .X(_0123_));
 sky130_fd_sc_hd__and3_1 _5223_ (.A(_0118_),
    .B(_0119_),
    .C(_0120_),
    .X(_0124_));
 sky130_fd_sc_hd__nand2_1 _5224_ (.A(net27),
    .B(net58),
    .Y(_0125_));
 sky130_fd_sc_hd__xnor2_1 _5225_ (.A(_4165_),
    .B(_4168_),
    .Y(_0126_));
 sky130_fd_sc_hd__xnor2_1 _5226_ (.A(_4203_),
    .B(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__or2_1 _5227_ (.A(_0125_),
    .B(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__a21o_1 _5228_ (.A1(_4174_),
    .A2(_4176_),
    .B1(_4201_),
    .X(_0129_));
 sky130_fd_sc_hd__or3_1 _5229_ (.A(_4173_),
    .B(_4175_),
    .C(_4202_),
    .X(_0130_));
 sky130_fd_sc_hd__nand4_2 _5230_ (.A(net26),
    .B(net58),
    .C(_0129_),
    .D(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__a22oi_1 _5231_ (.A1(net26),
    .A2(net58),
    .B1(_0129_),
    .B2(_0130_),
    .Y(_0133_));
 sky130_fd_sc_hd__a22o_1 _5232_ (.A1(net26),
    .A2(net58),
    .B1(_0129_),
    .B2(_0130_),
    .X(_0134_));
 sky130_fd_sc_hd__a2bb2o_1 _5233_ (.A1_N(_4180_),
    .A2_N(_4182_),
    .B1(_4188_),
    .B2(_4200_),
    .X(_0135_));
 sky130_fd_sc_hd__or4bb_1 _5234_ (.A(_4180_),
    .B(_4182_),
    .C_N(_4188_),
    .D_N(_4200_),
    .X(_0136_));
 sky130_fd_sc_hd__and4_1 _5235_ (.A(net23),
    .B(net58),
    .C(_0135_),
    .D(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__a22oi_1 _5236_ (.A1(net23),
    .A2(net58),
    .B1(_0135_),
    .B2(_0136_),
    .Y(_0138_));
 sky130_fd_sc_hd__a22o_1 _5237_ (.A1(net23),
    .A2(net58),
    .B1(_0135_),
    .B2(_0136_),
    .X(_0139_));
 sky130_fd_sc_hd__nand2_1 _5238_ (.A(net12),
    .B(net58),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _5239_ (.A(_0140_),
    .Y(_0141_));
 sky130_fd_sc_hd__xnor2_1 _5240_ (.A(_4183_),
    .B(_4186_),
    .Y(_0142_));
 sky130_fd_sc_hd__xnor2_2 _5241_ (.A(_4199_),
    .B(_0142_),
    .Y(_0144_));
 sky130_fd_sc_hd__and2_1 _5242_ (.A(_0141_),
    .B(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__nand2_1 _5243_ (.A(_0141_),
    .B(_0144_),
    .Y(_0146_));
 sky130_fd_sc_hd__a21oi_1 _5244_ (.A1(_4194_),
    .A2(_4195_),
    .B1(_4197_),
    .Y(_0147_));
 sky130_fd_sc_hd__a31o_1 _5245_ (.A1(_4194_),
    .A2(_4195_),
    .A3(_4197_),
    .B1(_0022_),
    .X(_0148_));
 sky130_fd_sc_hd__nor3_1 _5246_ (.A(_4198_),
    .B(_0147_),
    .C(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__o21a_1 _5247_ (.A1(_0141_),
    .A2(_0144_),
    .B1(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__o21ai_1 _5248_ (.A1(_0141_),
    .A2(_0144_),
    .B1(_0149_),
    .Y(_0151_));
 sky130_fd_sc_hd__o31ai_1 _5249_ (.A1(_0137_),
    .A2(_0145_),
    .A3(_0150_),
    .B1(_0139_),
    .Y(_0152_));
 sky130_fd_sc_hd__o31a_1 _5250_ (.A1(_0137_),
    .A2(_0145_),
    .A3(_0150_),
    .B1(_0139_),
    .X(_0153_));
 sky130_fd_sc_hd__a21o_1 _5251_ (.A1(_0131_),
    .A2(_0152_),
    .B1(_0133_),
    .X(_0155_));
 sky130_fd_sc_hd__a221o_1 _5252_ (.A1(_0125_),
    .A2(_0127_),
    .B1(_0131_),
    .B2(_0152_),
    .C1(_0133_),
    .X(_0156_));
 sky130_fd_sc_hd__a31o_1 _5253_ (.A1(_0123_),
    .A2(_0128_),
    .A3(_0156_),
    .B1(_0124_),
    .X(_0157_));
 sky130_fd_sc_hd__a31oi_1 _5254_ (.A1(_0123_),
    .A2(_0128_),
    .A3(_0156_),
    .B1(_0124_),
    .Y(_0158_));
 sky130_fd_sc_hd__a21o_1 _5255_ (.A1(_0115_),
    .A2(_0157_),
    .B1(_0116_),
    .X(_0159_));
 sky130_fd_sc_hd__o221a_1 _5256_ (.A1(_0106_),
    .A2(_0108_),
    .B1(_0114_),
    .B2(_0158_),
    .C1(_0117_),
    .X(_0160_));
 sky130_fd_sc_hd__o31a_1 _5257_ (.A1(_0104_),
    .A2(_0109_),
    .A3(_0160_),
    .B1(_0103_),
    .X(_0161_));
 sky130_fd_sc_hd__a21boi_2 _5258_ (.A1(_0096_),
    .A2(_0161_),
    .B1_N(_0097_),
    .Y(_0162_));
 sky130_fd_sc_hd__o21a_1 _5259_ (.A1(_0090_),
    .A2(_0162_),
    .B1(_0091_),
    .X(_0163_));
 sky130_fd_sc_hd__o211ai_2 _5260_ (.A1(_0090_),
    .A2(_0162_),
    .B1(_0091_),
    .C1(_0084_),
    .Y(_0164_));
 sky130_fd_sc_hd__a31o_1 _5261_ (.A1(_0076_),
    .A2(_0085_),
    .A3(_0164_),
    .B1(_0078_),
    .X(_0166_));
 sky130_fd_sc_hd__a21oi_1 _5262_ (.A1(_0071_),
    .A2(_0166_),
    .B1(_0072_),
    .Y(_0167_));
 sky130_fd_sc_hd__a211o_1 _5263_ (.A1(_0071_),
    .A2(_0166_),
    .B1(_0072_),
    .C1(_0065_),
    .X(_0168_));
 sky130_fd_sc_hd__a31o_1 _5264_ (.A1(_0060_),
    .A2(_0067_),
    .A3(_0168_),
    .B1(_0061_),
    .X(_0169_));
 sky130_fd_sc_hd__a311o_1 _5265_ (.A1(_0060_),
    .A2(_0067_),
    .A3(_0168_),
    .B1(_0061_),
    .C1(_0056_),
    .X(_0170_));
 sky130_fd_sc_hd__a31o_1 _5266_ (.A1(_0049_),
    .A2(_0054_),
    .A3(_0170_),
    .B1(_0047_),
    .X(_0171_));
 sky130_fd_sc_hd__a21oi_1 _5267_ (.A1(_0041_),
    .A2(_0171_),
    .B1(_0042_),
    .Y(_0172_));
 sky130_fd_sc_hd__a221o_1 _5268_ (.A1(_0035_),
    .A2(_0036_),
    .B1(_0041_),
    .B2(_0171_),
    .C1(_0042_),
    .X(_0173_));
 sky130_fd_sc_hd__nand2_1 _5269_ (.A(_0037_),
    .B(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__o211a_1 _5270_ (.A1(_0029_),
    .A2(_0031_),
    .B1(_0037_),
    .C1(_0173_),
    .X(_0175_));
 sky130_fd_sc_hd__o31ai_2 _5271_ (.A1(_0026_),
    .A2(_0032_),
    .A3(_0175_),
    .B1(_0025_),
    .Y(_0177_));
 sky130_fd_sc_hd__or2_1 _5272_ (.A(_0021_),
    .B(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_1 _5273_ (.A(net15),
    .B(net58),
    .Y(_0179_));
 sky130_fd_sc_hd__a21o_1 _5274_ (.A1(_0021_),
    .A2(_0177_),
    .B1(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__a21o_1 _5275_ (.A1(_0178_),
    .A2(_0180_),
    .B1(_0019_),
    .X(_0181_));
 sky130_fd_sc_hd__nand3_1 _5276_ (.A(_0019_),
    .B(_0178_),
    .C(_0180_),
    .Y(_0182_));
 sky130_fd_sc_hd__and3_1 _5277_ (.A(_3990_),
    .B(_0181_),
    .C(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__a21oi_1 _5278_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_3990_),
    .Y(_0184_));
 sky130_fd_sc_hd__a21o_1 _5279_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_3990_),
    .X(_0185_));
 sky130_fd_sc_hd__and2_1 _5280_ (.A(net13),
    .B(net59),
    .X(_0186_));
 sky130_fd_sc_hd__a211o_1 _5281_ (.A1(_0025_),
    .A2(_0027_),
    .B1(_0032_),
    .C1(_0175_),
    .X(_0188_));
 sky130_fd_sc_hd__o211ai_2 _5282_ (.A1(_0032_),
    .A2(_0175_),
    .B1(_0025_),
    .C1(_0027_),
    .Y(_0189_));
 sky130_fd_sc_hd__a21oi_1 _5283_ (.A1(_0188_),
    .A2(_0189_),
    .B1(_0186_),
    .Y(_0190_));
 sky130_fd_sc_hd__a21o_1 _5284_ (.A1(_0188_),
    .A2(_0189_),
    .B1(_0186_),
    .X(_0191_));
 sky130_fd_sc_hd__and3_1 _5285_ (.A(_0186_),
    .B(_0188_),
    .C(_0189_),
    .X(_0192_));
 sky130_fd_sc_hd__and2_1 _5286_ (.A(net11),
    .B(net59),
    .X(_0193_));
 sky130_fd_sc_hd__xnor2_1 _5287_ (.A(_0028_),
    .B(_0031_),
    .Y(_0194_));
 sky130_fd_sc_hd__xnor2_1 _5288_ (.A(_0174_),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__or2_1 _5289_ (.A(_0193_),
    .B(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__nand2_1 _5290_ (.A(net10),
    .B(net59),
    .Y(_0197_));
 sky130_fd_sc_hd__xor2_1 _5291_ (.A(_0035_),
    .B(_0036_),
    .X(_0199_));
 sky130_fd_sc_hd__xnor2_1 _5292_ (.A(_0172_),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__a21o_1 _5293_ (.A1(net10),
    .A2(net59),
    .B1(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__and3_1 _5294_ (.A(net10),
    .B(net59),
    .C(_0200_),
    .X(_0202_));
 sky130_fd_sc_hd__a21o_1 _5295_ (.A1(_0041_),
    .A2(_0043_),
    .B1(_0171_),
    .X(_0203_));
 sky130_fd_sc_hd__nand3_1 _5296_ (.A(_0041_),
    .B(_0043_),
    .C(_0171_),
    .Y(_0204_));
 sky130_fd_sc_hd__and4_1 _5297_ (.A(net9),
    .B(net59),
    .C(_0203_),
    .D(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__a22oi_2 _5298_ (.A1(net9),
    .A2(net59),
    .B1(_0203_),
    .B2(_0204_),
    .Y(_0206_));
 sky130_fd_sc_hd__a22o_1 _5299_ (.A1(net9),
    .A2(net59),
    .B1(_0203_),
    .B2(_0204_),
    .X(_0207_));
 sky130_fd_sc_hd__nand2_1 _5300_ (.A(net8),
    .B(net59),
    .Y(_0208_));
 sky130_fd_sc_hd__o211ai_2 _5301_ (.A1(_0047_),
    .A2(_0048_),
    .B1(_0054_),
    .C1(_0170_),
    .Y(_0210_));
 sky130_fd_sc_hd__a211o_1 _5302_ (.A1(_0054_),
    .A2(_0170_),
    .B1(_0047_),
    .C1(_0048_),
    .X(_0211_));
 sky130_fd_sc_hd__a21oi_1 _5303_ (.A1(_0210_),
    .A2(_0211_),
    .B1(_0208_),
    .Y(_0212_));
 sky130_fd_sc_hd__and3_1 _5304_ (.A(_0208_),
    .B(_0210_),
    .C(_0211_),
    .X(_0213_));
 sky130_fd_sc_hd__nand3_1 _5305_ (.A(_0208_),
    .B(_0210_),
    .C(_0211_),
    .Y(_0214_));
 sky130_fd_sc_hd__nand2_1 _5306_ (.A(net7),
    .B(net59),
    .Y(_0215_));
 sky130_fd_sc_hd__nor2_1 _5307_ (.A(_0053_),
    .B(_0056_),
    .Y(_0216_));
 sky130_fd_sc_hd__xor2_1 _5308_ (.A(_0169_),
    .B(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__nand2b_1 _5309_ (.A_N(_0217_),
    .B(_0215_),
    .Y(_0218_));
 sky130_fd_sc_hd__and3_1 _5310_ (.A(net7),
    .B(net59),
    .C(_0217_),
    .X(_0219_));
 sky130_fd_sc_hd__xnor2_1 _5311_ (.A(_0057_),
    .B(_0059_),
    .Y(_0221_));
 sky130_fd_sc_hd__a21o_1 _5312_ (.A1(_0067_),
    .A2(_0168_),
    .B1(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__nand3_1 _5313_ (.A(_0067_),
    .B(_0168_),
    .C(_0221_),
    .Y(_0223_));
 sky130_fd_sc_hd__a22oi_2 _5314_ (.A1(net6),
    .A2(net59),
    .B1(_0222_),
    .B2(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_2 _5315_ (.A(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__nand4_2 _5316_ (.A(net6),
    .B(net59),
    .C(_0222_),
    .D(_0223_),
    .Y(_0226_));
 sky130_fd_sc_hd__and2_1 _5317_ (.A(net5),
    .B(net59),
    .X(_0227_));
 sky130_fd_sc_hd__and2b_1 _5318_ (.A_N(_0065_),
    .B(_0067_),
    .X(_0228_));
 sky130_fd_sc_hd__xnor2_2 _5319_ (.A(_0167_),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__nand2_1 _5320_ (.A(_0227_),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _5321_ (.A(net4),
    .B(net59),
    .Y(_0232_));
 sky130_fd_sc_hd__xnor2_1 _5322_ (.A(_0068_),
    .B(_0070_),
    .Y(_0233_));
 sky130_fd_sc_hd__xnor2_1 _5323_ (.A(_0166_),
    .B(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__and3_1 _5324_ (.A(net4),
    .B(net59),
    .C(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__nand2b_1 _5325_ (.A_N(_0234_),
    .B(_0232_),
    .Y(_0236_));
 sky130_fd_sc_hd__xnor2_1 _5326_ (.A(_0073_),
    .B(_0075_),
    .Y(_0237_));
 sky130_fd_sc_hd__a21o_1 _5327_ (.A1(_0085_),
    .A2(_0164_),
    .B1(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__nand3_1 _5328_ (.A(_0085_),
    .B(_0164_),
    .C(_0237_),
    .Y(_0239_));
 sky130_fd_sc_hd__and4_1 _5329_ (.A(net3),
    .B(net59),
    .C(_0238_),
    .D(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__nand4_1 _5330_ (.A(net3),
    .B(net59),
    .C(_0238_),
    .D(_0239_),
    .Y(_0241_));
 sky130_fd_sc_hd__a22o_1 _5331_ (.A1(net3),
    .A2(net59),
    .B1(_0238_),
    .B2(_0239_),
    .X(_0243_));
 sky130_fd_sc_hd__nand2_1 _5332_ (.A(net2),
    .B(net59),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_2 _5333_ (.A(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__xor2_1 _5334_ (.A(_0079_),
    .B(_0083_),
    .X(_0246_));
 sky130_fd_sc_hd__xnor2_1 _5335_ (.A(_0163_),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__and2_1 _5336_ (.A(_0245_),
    .B(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__nand2_1 _5337_ (.A(net32),
    .B(net59),
    .Y(_0249_));
 sky130_fd_sc_hd__xnor2_1 _5338_ (.A(_0086_),
    .B(_0089_),
    .Y(_0250_));
 sky130_fd_sc_hd__xnor2_1 _5339_ (.A(_0162_),
    .B(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__and3_1 _5340_ (.A(net32),
    .B(net59),
    .C(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__a21o_1 _5341_ (.A1(net32),
    .A2(net59),
    .B1(_0251_),
    .X(_0254_));
 sky130_fd_sc_hd__a21o_1 _5342_ (.A1(_0096_),
    .A2(_0097_),
    .B1(_0161_),
    .X(_0255_));
 sky130_fd_sc_hd__nand3_1 _5343_ (.A(_0096_),
    .B(_0097_),
    .C(_0161_),
    .Y(_0256_));
 sky130_fd_sc_hd__and4_1 _5344_ (.A(net31),
    .B(net59),
    .C(_0255_),
    .D(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__a22oi_1 _5345_ (.A1(net31),
    .A2(net59),
    .B1(_0255_),
    .B2(_0256_),
    .Y(_0258_));
 sky130_fd_sc_hd__a22o_1 _5346_ (.A1(net31),
    .A2(net59),
    .B1(_0255_),
    .B2(_0256_),
    .X(_0259_));
 sky130_fd_sc_hd__and2_1 _5347_ (.A(net30),
    .B(net59),
    .X(_0260_));
 sky130_fd_sc_hd__o22a_1 _5348_ (.A1(_0102_),
    .A2(_0104_),
    .B1(_0109_),
    .B2(_0160_),
    .X(_0261_));
 sky130_fd_sc_hd__or4_1 _5349_ (.A(_0102_),
    .B(_0104_),
    .C(_0109_),
    .D(_0160_),
    .X(_0262_));
 sky130_fd_sc_hd__nand2b_1 _5350_ (.A_N(_0261_),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__or2_1 _5351_ (.A(_0260_),
    .B(_0263_),
    .X(_0265_));
 sky130_fd_sc_hd__nand2_1 _5352_ (.A(net29),
    .B(net59),
    .Y(_0266_));
 sky130_fd_sc_hd__xnor2_1 _5353_ (.A(_0105_),
    .B(_0108_),
    .Y(_0267_));
 sky130_fd_sc_hd__xnor2_1 _5354_ (.A(_0159_),
    .B(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__a21o_1 _5355_ (.A1(net29),
    .A2(net59),
    .B1(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__and3_1 _5356_ (.A(net29),
    .B(net59),
    .C(_0268_),
    .X(_0270_));
 sky130_fd_sc_hd__nand2_1 _5357_ (.A(net28),
    .B(net59),
    .Y(_0271_));
 sky130_fd_sc_hd__a21o_1 _5358_ (.A1(_0115_),
    .A2(_0117_),
    .B1(_0157_),
    .X(_0272_));
 sky130_fd_sc_hd__or3_1 _5359_ (.A(_0114_),
    .B(_0116_),
    .C(_0158_),
    .X(_0273_));
 sky130_fd_sc_hd__nand3_1 _5360_ (.A(_0271_),
    .B(_0272_),
    .C(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__a21o_1 _5361_ (.A1(_0272_),
    .A2(_0273_),
    .B1(_0271_),
    .X(_0276_));
 sky130_fd_sc_hd__nand2_1 _5362_ (.A(net27),
    .B(net59),
    .Y(_0277_));
 sky130_fd_sc_hd__a2bb2o_1 _5363_ (.A1_N(_0122_),
    .A2_N(_0124_),
    .B1(_0128_),
    .B2(_0156_),
    .X(_0278_));
 sky130_fd_sc_hd__or4bb_1 _5364_ (.A(_0122_),
    .B(_0124_),
    .C_N(_0128_),
    .D_N(_0156_),
    .X(_0279_));
 sky130_fd_sc_hd__a21oi_1 _5365_ (.A1(_0278_),
    .A2(_0279_),
    .B1(_0277_),
    .Y(_0280_));
 sky130_fd_sc_hd__a21o_1 _5366_ (.A1(_0278_),
    .A2(_0279_),
    .B1(_0277_),
    .X(_0281_));
 sky130_fd_sc_hd__and3_1 _5367_ (.A(_0277_),
    .B(_0278_),
    .C(_0279_),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _5368_ (.A(net26),
    .B(net59),
    .Y(_0283_));
 sky130_fd_sc_hd__xnor2_1 _5369_ (.A(_0125_),
    .B(_0127_),
    .Y(_0284_));
 sky130_fd_sc_hd__xnor2_1 _5370_ (.A(_0155_),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__or2_1 _5371_ (.A(_0283_),
    .B(_0285_),
    .X(_0287_));
 sky130_fd_sc_hd__a21o_1 _5372_ (.A1(_0131_),
    .A2(_0134_),
    .B1(_0153_),
    .X(_0288_));
 sky130_fd_sc_hd__nand3_1 _5373_ (.A(_0131_),
    .B(_0134_),
    .C(_0153_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand4_2 _5374_ (.A(net23),
    .B(net59),
    .C(_0288_),
    .D(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__a22oi_1 _5375_ (.A1(net23),
    .A2(net59),
    .B1(_0288_),
    .B2(_0289_),
    .Y(_0291_));
 sky130_fd_sc_hd__a22o_1 _5376_ (.A1(net23),
    .A2(net59),
    .B1(_0288_),
    .B2(_0289_),
    .X(_0292_));
 sky130_fd_sc_hd__o211ai_1 _5377_ (.A1(_0137_),
    .A2(_0138_),
    .B1(_0146_),
    .C1(_0151_),
    .Y(_0293_));
 sky130_fd_sc_hd__a211o_1 _5378_ (.A1(_0146_),
    .A2(_0151_),
    .B1(_0137_),
    .C1(_0138_),
    .X(_0294_));
 sky130_fd_sc_hd__nand4_1 _5379_ (.A(net12),
    .B(net59),
    .C(_0293_),
    .D(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__a22o_1 _5380_ (.A1(net12),
    .A2(net59),
    .B1(_0293_),
    .B2(_0294_),
    .X(_0296_));
 sky130_fd_sc_hd__xnor2_1 _5381_ (.A(_0140_),
    .B(_0144_),
    .Y(_0298_));
 sky130_fd_sc_hd__a21oi_1 _5382_ (.A1(_0149_),
    .A2(_0298_),
    .B1(_4198_),
    .Y(_0299_));
 sky130_fd_sc_hd__o211a_1 _5383_ (.A1(_0149_),
    .A2(_0298_),
    .B1(_0299_),
    .C1(net59),
    .X(_0300_));
 sky130_fd_sc_hd__a21boi_2 _5384_ (.A1(_0296_),
    .A2(_0300_),
    .B1_N(_0295_),
    .Y(_0301_));
 sky130_fd_sc_hd__a21oi_1 _5385_ (.A1(_0290_),
    .A2(_0301_),
    .B1(_0291_),
    .Y(_0302_));
 sky130_fd_sc_hd__a221o_1 _5386_ (.A1(_0283_),
    .A2(_0285_),
    .B1(_0290_),
    .B2(_0301_),
    .C1(_0291_),
    .X(_0303_));
 sky130_fd_sc_hd__a31oi_2 _5387_ (.A1(_0281_),
    .A2(_0287_),
    .A3(_0303_),
    .B1(_0282_),
    .Y(_0304_));
 sky130_fd_sc_hd__a21bo_1 _5388_ (.A1(_0274_),
    .A2(_0304_),
    .B1_N(_0276_),
    .X(_0305_));
 sky130_fd_sc_hd__a21oi_1 _5389_ (.A1(_0269_),
    .A2(_0305_),
    .B1(_0270_),
    .Y(_0306_));
 sky130_fd_sc_hd__a221o_1 _5390_ (.A1(_0260_),
    .A2(_0263_),
    .B1(_0269_),
    .B2(_0305_),
    .C1(_0270_),
    .X(_0307_));
 sky130_fd_sc_hd__a31o_1 _5391_ (.A1(_0259_),
    .A2(_0265_),
    .A3(_0307_),
    .B1(_0257_),
    .X(_0309_));
 sky130_fd_sc_hd__o21a_1 _5392_ (.A1(_0252_),
    .A2(_0309_),
    .B1(_0254_),
    .X(_0310_));
 sky130_fd_sc_hd__o221a_1 _5393_ (.A1(_0245_),
    .A2(_0247_),
    .B1(_0252_),
    .B2(_0309_),
    .C1(_0254_),
    .X(_0311_));
 sky130_fd_sc_hd__o31a_2 _5394_ (.A1(_0240_),
    .A2(_0248_),
    .A3(_0311_),
    .B1(_0243_),
    .X(_0312_));
 sky130_fd_sc_hd__o21ai_1 _5395_ (.A1(_0235_),
    .A2(_0312_),
    .B1(_0236_),
    .Y(_0313_));
 sky130_fd_sc_hd__o221ai_4 _5396_ (.A1(_0227_),
    .A2(_0229_),
    .B1(_0235_),
    .B2(_0312_),
    .C1(_0236_),
    .Y(_0314_));
 sky130_fd_sc_hd__nand2_1 _5397_ (.A(_0230_),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand3_1 _5398_ (.A(_0226_),
    .B(_0230_),
    .C(_0314_),
    .Y(_0316_));
 sky130_fd_sc_hd__a21o_1 _5399_ (.A1(_0230_),
    .A2(_0314_),
    .B1(_0224_),
    .X(_0317_));
 sky130_fd_sc_hd__a31oi_1 _5400_ (.A1(_0218_),
    .A2(_0225_),
    .A3(_0316_),
    .B1(_0219_),
    .Y(_0318_));
 sky130_fd_sc_hd__a311o_1 _5401_ (.A1(_0218_),
    .A2(_0225_),
    .A3(_0316_),
    .B1(_0219_),
    .C1(_0212_),
    .X(_0320_));
 sky130_fd_sc_hd__a31o_1 _5402_ (.A1(_0207_),
    .A2(_0214_),
    .A3(_0320_),
    .B1(_0205_),
    .X(_0321_));
 sky130_fd_sc_hd__a21o_1 _5403_ (.A1(_0201_),
    .A2(_0321_),
    .B1(_0202_),
    .X(_0322_));
 sky130_fd_sc_hd__a221o_1 _5404_ (.A1(_0193_),
    .A2(_0195_),
    .B1(_0201_),
    .B2(_0321_),
    .C1(_0202_),
    .X(_0323_));
 sky130_fd_sc_hd__nand2_1 _5405_ (.A(_0196_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__a31o_1 _5406_ (.A1(_0191_),
    .A2(_0196_),
    .A3(_0323_),
    .B1(_0192_),
    .X(_0325_));
 sky130_fd_sc_hd__xor2_1 _5407_ (.A(_0021_),
    .B(_0177_),
    .X(_0326_));
 sky130_fd_sc_hd__xnor2_1 _5408_ (.A(_0179_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__nor2_1 _5409_ (.A(_0325_),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__and2_1 _5410_ (.A(net14),
    .B(net59),
    .X(_0329_));
 sky130_fd_sc_hd__a21oi_1 _5411_ (.A1(_0325_),
    .A2(_0327_),
    .B1(_0329_),
    .Y(_0331_));
 sky130_fd_sc_hd__nor3_1 _5412_ (.A(_0183_),
    .B(_0328_),
    .C(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__o31a_1 _5413_ (.A1(_0183_),
    .A2(_0328_),
    .A3(_0331_),
    .B1(_0185_),
    .X(_0333_));
 sky130_fd_sc_hd__a2bb2oi_1 _5414_ (.A1_N(_0017_),
    .A2_N(_0018_),
    .B1(_0178_),
    .B2(_0180_),
    .Y(_0334_));
 sky130_fd_sc_hd__a21o_1 _5415_ (.A1(net58),
    .A2(_0017_),
    .B1(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__o311a_1 _5416_ (.A1(_0184_),
    .A2(_0332_),
    .A3(_0335_),
    .B1(_1716_),
    .C1(net59),
    .X(_0336_));
 sky130_fd_sc_hd__a21o_1 _5417_ (.A1(net60),
    .A2(_1716_),
    .B1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__a21bo_1 _5418_ (.A1(net60),
    .A2(_0336_),
    .B1_N(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__o22ai_1 _5419_ (.A1(_0183_),
    .A2(_0184_),
    .B1(_0328_),
    .B2(_0331_),
    .Y(_0339_));
 sky130_fd_sc_hd__or4_1 _5420_ (.A(_0183_),
    .B(_0184_),
    .C(_0328_),
    .D(_0331_),
    .X(_0340_));
 sky130_fd_sc_hd__and4_1 _5421_ (.A(net14),
    .B(net60),
    .C(_0339_),
    .D(_0340_),
    .X(_0342_));
 sky130_fd_sc_hd__a22o_1 _5422_ (.A1(net14),
    .A2(net60),
    .B1(_0339_),
    .B2(_0340_),
    .X(_0343_));
 sky130_fd_sc_hd__xor2_1 _5423_ (.A(_0325_),
    .B(_0327_),
    .X(_0344_));
 sky130_fd_sc_hd__xnor2_1 _5424_ (.A(_0329_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__and2_1 _5425_ (.A(net11),
    .B(net60),
    .X(_0346_));
 sky130_fd_sc_hd__or2_1 _5426_ (.A(_0190_),
    .B(_0192_),
    .X(_0347_));
 sky130_fd_sc_hd__xor2_2 _5427_ (.A(_0324_),
    .B(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__nand2_1 _5428_ (.A(_0346_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__nand2_1 _5429_ (.A(net10),
    .B(net60),
    .Y(_0350_));
 sky130_fd_sc_hd__xnor2_1 _5430_ (.A(_0193_),
    .B(_0195_),
    .Y(_0351_));
 sky130_fd_sc_hd__xnor2_1 _5431_ (.A(_0322_),
    .B(_0351_),
    .Y(_0353_));
 sky130_fd_sc_hd__a21o_1 _5432_ (.A1(net10),
    .A2(net60),
    .B1(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__and3_1 _5433_ (.A(net10),
    .B(net60),
    .C(_0353_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _5434_ (.A(net9),
    .B(net60),
    .X(_0356_));
 sky130_fd_sc_hd__xor2_1 _5435_ (.A(_0197_),
    .B(_0200_),
    .X(_0357_));
 sky130_fd_sc_hd__xnor2_1 _5436_ (.A(_0321_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__and2_1 _5437_ (.A(_0356_),
    .B(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__nor2_1 _5438_ (.A(_0356_),
    .B(_0358_),
    .Y(_0360_));
 sky130_fd_sc_hd__or2_1 _5439_ (.A(_0356_),
    .B(_0358_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_1 _5440_ (.A(net8),
    .B(net60),
    .Y(_0362_));
 sky130_fd_sc_hd__o211ai_2 _5441_ (.A1(_0205_),
    .A2(_0206_),
    .B1(_0214_),
    .C1(_0320_),
    .Y(_0364_));
 sky130_fd_sc_hd__a211o_1 _5442_ (.A1(_0214_),
    .A2(_0320_),
    .B1(_0205_),
    .C1(_0206_),
    .X(_0365_));
 sky130_fd_sc_hd__and3_1 _5443_ (.A(_0362_),
    .B(_0364_),
    .C(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__nand3_1 _5444_ (.A(_0362_),
    .B(_0364_),
    .C(_0365_),
    .Y(_0367_));
 sky130_fd_sc_hd__a21oi_1 _5445_ (.A1(_0364_),
    .A2(_0365_),
    .B1(_0362_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_1 _5446_ (.A(net7),
    .B(net60),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _5447_ (.A(_0212_),
    .B(_0213_),
    .Y(_0370_));
 sky130_fd_sc_hd__xnor2_1 _5448_ (.A(_0318_),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__and3_1 _5449_ (.A(net7),
    .B(net60),
    .C(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__a21o_1 _5450_ (.A1(net7),
    .A2(net60),
    .B1(_0371_),
    .X(_0373_));
 sky130_fd_sc_hd__xor2_1 _5451_ (.A(_0215_),
    .B(_0217_),
    .X(_0375_));
 sky130_fd_sc_hd__nand3_1 _5452_ (.A(_0226_),
    .B(_0317_),
    .C(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__a21o_1 _5453_ (.A1(_0226_),
    .A2(_0317_),
    .B1(_0375_),
    .X(_0377_));
 sky130_fd_sc_hd__a22o_1 _5454_ (.A1(net6),
    .A2(net60),
    .B1(_0376_),
    .B2(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__nand4_2 _5455_ (.A(net6),
    .B(net60),
    .C(_0376_),
    .D(_0377_),
    .Y(_0379_));
 sky130_fd_sc_hd__and2_1 _5456_ (.A(net5),
    .B(net60),
    .X(_0380_));
 sky130_fd_sc_hd__nand2b_1 _5457_ (.A_N(_0224_),
    .B(_0226_),
    .Y(_0381_));
 sky130_fd_sc_hd__xnor2_2 _5458_ (.A(_0315_),
    .B(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_1 _5459_ (.A(_0380_),
    .B(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand2_1 _5460_ (.A(net4),
    .B(net60),
    .Y(_0384_));
 sky130_fd_sc_hd__xor2_1 _5461_ (.A(_0227_),
    .B(_0229_),
    .X(_0386_));
 sky130_fd_sc_hd__xnor2_1 _5462_ (.A(_0313_),
    .B(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__and3_1 _5463_ (.A(net4),
    .B(net60),
    .C(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__a21o_1 _5464_ (.A1(net4),
    .A2(net60),
    .B1(_0387_),
    .X(_0389_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(net3),
    .B(net60),
    .Y(_0390_));
 sky130_fd_sc_hd__xor2_1 _5466_ (.A(_0232_),
    .B(_0234_),
    .X(_0391_));
 sky130_fd_sc_hd__xnor2_1 _5467_ (.A(_0312_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__a21o_1 _5468_ (.A1(net3),
    .A2(net60),
    .B1(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__and3_1 _5469_ (.A(net3),
    .B(net60),
    .C(_0392_),
    .X(_0394_));
 sky130_fd_sc_hd__nand2_1 _5470_ (.A(net2),
    .B(net60),
    .Y(_0395_));
 sky130_fd_sc_hd__inv_2 _5471_ (.A(_0395_),
    .Y(_0397_));
 sky130_fd_sc_hd__a211o_1 _5472_ (.A1(_0241_),
    .A2(_0243_),
    .B1(_0248_),
    .C1(_0311_),
    .X(_0398_));
 sky130_fd_sc_hd__o211ai_1 _5473_ (.A1(_0248_),
    .A2(_0311_),
    .B1(_0241_),
    .C1(_0243_),
    .Y(_0399_));
 sky130_fd_sc_hd__and3_1 _5474_ (.A(_0397_),
    .B(_0398_),
    .C(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__a21o_1 _5475_ (.A1(_0398_),
    .A2(_0399_),
    .B1(_0397_),
    .X(_0401_));
 sky130_fd_sc_hd__nand2_1 _5476_ (.A(net32),
    .B(net60),
    .Y(_0402_));
 sky130_fd_sc_hd__xnor2_1 _5477_ (.A(_0245_),
    .B(_0247_),
    .Y(_0403_));
 sky130_fd_sc_hd__xnor2_1 _5478_ (.A(_0310_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__and3_1 _5479_ (.A(net32),
    .B(net60),
    .C(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__nand2b_1 _5480_ (.A_N(_0404_),
    .B(_0402_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_1 _5481_ (.A(net31),
    .B(net60),
    .Y(_0408_));
 sky130_fd_sc_hd__xor2_1 _5482_ (.A(_0249_),
    .B(_0251_),
    .X(_0409_));
 sky130_fd_sc_hd__xnor2_1 _5483_ (.A(_0309_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2b_1 _5484_ (.A_N(_0410_),
    .B(_0408_),
    .Y(_0411_));
 sky130_fd_sc_hd__and3_1 _5485_ (.A(net31),
    .B(net60),
    .C(_0410_),
    .X(_0412_));
 sky130_fd_sc_hd__a2bb2o_1 _5486_ (.A1_N(_0257_),
    .A2_N(_0258_),
    .B1(_0265_),
    .B2(_0307_),
    .X(_0413_));
 sky130_fd_sc_hd__or4bb_1 _5487_ (.A(_0257_),
    .B(_0258_),
    .C_N(_0265_),
    .D_N(_0307_),
    .X(_0414_));
 sky130_fd_sc_hd__and4_1 _5488_ (.A(net30),
    .B(net60),
    .C(_0413_),
    .D(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__a22oi_1 _5489_ (.A1(net30),
    .A2(net60),
    .B1(_0413_),
    .B2(_0414_),
    .Y(_0416_));
 sky130_fd_sc_hd__a22o_1 _5490_ (.A1(net30),
    .A2(net60),
    .B1(_0413_),
    .B2(_0414_),
    .X(_0417_));
 sky130_fd_sc_hd__and2_1 _5491_ (.A(net29),
    .B(net60),
    .X(_0419_));
 sky130_fd_sc_hd__xor2_1 _5492_ (.A(_0260_),
    .B(_0263_),
    .X(_0420_));
 sky130_fd_sc_hd__xnor2_1 _5493_ (.A(_0306_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__and2_1 _5494_ (.A(_0419_),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_1 _5495_ (.A(net28),
    .B(net60),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_2 _5496_ (.A(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__xor2_1 _5497_ (.A(_0266_),
    .B(_0268_),
    .X(_0425_));
 sky130_fd_sc_hd__xnor2_1 _5498_ (.A(_0305_),
    .B(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__and2_1 _5499_ (.A(_0424_),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__a21o_1 _5500_ (.A1(_0274_),
    .A2(_0276_),
    .B1(_0304_),
    .X(_0428_));
 sky130_fd_sc_hd__nand3_1 _5501_ (.A(_0274_),
    .B(_0276_),
    .C(_0304_),
    .Y(_0430_));
 sky130_fd_sc_hd__and4_1 _5502_ (.A(net27),
    .B(net60),
    .C(_0428_),
    .D(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__o2bb2a_1 _5503_ (.A1_N(_0428_),
    .A2_N(_0430_),
    .B1(_4187_),
    .B2(_0033_),
    .X(_0432_));
 sky130_fd_sc_hd__a22o_1 _5504_ (.A1(net27),
    .A2(net60),
    .B1(_0428_),
    .B2(_0430_),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _5505_ (.A(net26),
    .B(net60),
    .X(_0434_));
 sky130_fd_sc_hd__o211ai_2 _5506_ (.A1(_0280_),
    .A2(_0282_),
    .B1(_0287_),
    .C1(_0303_),
    .Y(_0435_));
 sky130_fd_sc_hd__a211o_1 _5507_ (.A1(_0287_),
    .A2(_0303_),
    .B1(_0280_),
    .C1(_0282_),
    .X(_0436_));
 sky130_fd_sc_hd__a21oi_1 _5508_ (.A1(_0435_),
    .A2(_0436_),
    .B1(_0434_),
    .Y(_0437_));
 sky130_fd_sc_hd__a21o_1 _5509_ (.A1(_0435_),
    .A2(_0436_),
    .B1(_0434_),
    .X(_0438_));
 sky130_fd_sc_hd__and3_1 _5510_ (.A(_0434_),
    .B(_0435_),
    .C(_0436_),
    .X(_0439_));
 sky130_fd_sc_hd__nand2_1 _5511_ (.A(net23),
    .B(net60),
    .Y(_0441_));
 sky130_fd_sc_hd__xnor2_1 _5512_ (.A(_0283_),
    .B(_0285_),
    .Y(_0442_));
 sky130_fd_sc_hd__xnor2_1 _5513_ (.A(_0302_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand2b_1 _5514_ (.A_N(_0443_),
    .B(_0441_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _5515_ (.A(net12),
    .B(net60),
    .Y(_0445_));
 sky130_fd_sc_hd__nand3_1 _5516_ (.A(_0290_),
    .B(_0292_),
    .C(_0301_),
    .Y(_0446_));
 sky130_fd_sc_hd__a21o_1 _5517_ (.A1(_0290_),
    .A2(_0292_),
    .B1(_0301_),
    .X(_0447_));
 sky130_fd_sc_hd__a21oi_1 _5518_ (.A1(_0446_),
    .A2(_0447_),
    .B1(_0445_),
    .Y(_0448_));
 sky130_fd_sc_hd__and3_1 _5519_ (.A(_0445_),
    .B(_0446_),
    .C(_0447_),
    .X(_0449_));
 sky130_fd_sc_hd__a21oi_1 _5520_ (.A1(_0295_),
    .A2(_0296_),
    .B1(_0300_),
    .Y(_0450_));
 sky130_fd_sc_hd__a31o_1 _5521_ (.A1(_0295_),
    .A2(_0296_),
    .A3(_0300_),
    .B1(_0033_),
    .X(_0452_));
 sky130_fd_sc_hd__nor3_1 _5522_ (.A(_4198_),
    .B(_0450_),
    .C(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__or3_1 _5523_ (.A(_4198_),
    .B(_0450_),
    .C(_0452_),
    .X(_0454_));
 sky130_fd_sc_hd__a31oi_1 _5524_ (.A1(_0445_),
    .A2(_0446_),
    .A3(_0447_),
    .B1(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__nor2_1 _5525_ (.A(_0448_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__a311o_1 _5526_ (.A1(net23),
    .A2(net60),
    .A3(_0443_),
    .B1(_0448_),
    .C1(_0455_),
    .X(_0457_));
 sky130_fd_sc_hd__a31o_1 _5527_ (.A1(_0438_),
    .A2(_0444_),
    .A3(_0457_),
    .B1(_0439_),
    .X(_0458_));
 sky130_fd_sc_hd__o21ai_1 _5528_ (.A1(_0431_),
    .A2(_0458_),
    .B1(_0433_),
    .Y(_0459_));
 sky130_fd_sc_hd__o221a_1 _5529_ (.A1(_0424_),
    .A2(_0426_),
    .B1(_0431_),
    .B2(_0458_),
    .C1(_0433_),
    .X(_0460_));
 sky130_fd_sc_hd__or2_1 _5530_ (.A(_0427_),
    .B(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__o22a_1 _5531_ (.A1(_0419_),
    .A2(_0421_),
    .B1(_0427_),
    .B2(_0460_),
    .X(_0463_));
 sky130_fd_sc_hd__o31a_1 _5532_ (.A1(_0415_),
    .A2(_0422_),
    .A3(_0463_),
    .B1(_0417_),
    .X(_0464_));
 sky130_fd_sc_hd__or2_1 _5533_ (.A(_0412_),
    .B(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__a21o_1 _5534_ (.A1(_0411_),
    .A2(_0464_),
    .B1(_0412_),
    .X(_0466_));
 sky130_fd_sc_hd__o21ai_1 _5535_ (.A1(_0405_),
    .A2(_0466_),
    .B1(_0406_),
    .Y(_0467_));
 sky130_fd_sc_hd__a311o_1 _5536_ (.A1(_0406_),
    .A2(_0411_),
    .A3(_0465_),
    .B1(_0405_),
    .C1(_0400_),
    .X(_0468_));
 sky130_fd_sc_hd__a31o_2 _5537_ (.A1(_0393_),
    .A2(_0401_),
    .A3(_0468_),
    .B1(_0394_),
    .X(_0469_));
 sky130_fd_sc_hd__o21ai_1 _5538_ (.A1(_0388_),
    .A2(_0469_),
    .B1(_0389_),
    .Y(_0470_));
 sky130_fd_sc_hd__o221ai_4 _5539_ (.A1(_0380_),
    .A2(_0382_),
    .B1(_0388_),
    .B2(_0469_),
    .C1(_0389_),
    .Y(_0471_));
 sky130_fd_sc_hd__nand3_1 _5540_ (.A(_0379_),
    .B(_0383_),
    .C(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__a21bo_1 _5541_ (.A1(_0383_),
    .A2(_0471_),
    .B1_N(_0378_),
    .X(_0474_));
 sky130_fd_sc_hd__a31o_1 _5542_ (.A1(_0373_),
    .A2(_0378_),
    .A3(_0472_),
    .B1(_0372_),
    .X(_0475_));
 sky130_fd_sc_hd__a311o_1 _5543_ (.A1(_0373_),
    .A2(_0378_),
    .A3(_0472_),
    .B1(_0372_),
    .C1(_0368_),
    .X(_0476_));
 sky130_fd_sc_hd__a31o_1 _5544_ (.A1(_0361_),
    .A2(_0367_),
    .A3(_0476_),
    .B1(_0359_),
    .X(_0477_));
 sky130_fd_sc_hd__o21ai_1 _5545_ (.A1(_0355_),
    .A2(_0477_),
    .B1(_0354_),
    .Y(_0478_));
 sky130_fd_sc_hd__o221ai_4 _5546_ (.A1(_0346_),
    .A2(_0348_),
    .B1(_0355_),
    .B2(_0477_),
    .C1(_0354_),
    .Y(_0479_));
 sky130_fd_sc_hd__nand3_1 _5547_ (.A(_0345_),
    .B(_0349_),
    .C(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a21oi_1 _5548_ (.A1(_0349_),
    .A2(_0479_),
    .B1(_0345_),
    .Y(_0481_));
 sky130_fd_sc_hd__a21o_1 _5549_ (.A1(_0349_),
    .A2(_0479_),
    .B1(_0345_),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _5550_ (.A(net13),
    .B(net60),
    .Y(_0483_));
 sky130_fd_sc_hd__a311oi_1 _5551_ (.A1(_0345_),
    .A2(_0349_),
    .A3(_0479_),
    .B1(_0033_),
    .C1(_0000_),
    .Y(_0485_));
 sky130_fd_sc_hd__or2_1 _5552_ (.A(_0481_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__o31a_1 _5553_ (.A1(_0342_),
    .A2(_0481_),
    .A3(_0485_),
    .B1(_0343_),
    .X(_0487_));
 sky130_fd_sc_hd__xnor2_1 _5554_ (.A(_0333_),
    .B(_0335_),
    .Y(_0488_));
 sky130_fd_sc_hd__xnor2_1 _5555_ (.A(_3989_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__nor2_1 _5556_ (.A(_0487_),
    .B(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__nand2_1 _5557_ (.A(_0487_),
    .B(_0489_),
    .Y(_0491_));
 sky130_fd_sc_hd__nand2_1 _5558_ (.A(net15),
    .B(net60),
    .Y(_0492_));
 sky130_fd_sc_hd__o21ai_1 _5559_ (.A1(_0490_),
    .A2(_0492_),
    .B1(_0491_),
    .Y(_0493_));
 sky130_fd_sc_hd__xnor2_1 _5560_ (.A(_0338_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__and3_1 _5561_ (.A(net15),
    .B(net61),
    .C(_0494_),
    .X(_0496_));
 sky130_fd_sc_hd__a21o_1 _5562_ (.A1(net15),
    .A2(net61),
    .B1(_0494_),
    .X(_0497_));
 sky130_fd_sc_hd__nand2_1 _5563_ (.A(net13),
    .B(net61),
    .Y(_0498_));
 sky130_fd_sc_hd__nand2b_1 _5564_ (.A_N(_0342_),
    .B(_0343_),
    .Y(_0499_));
 sky130_fd_sc_hd__xnor2_1 _5565_ (.A(_0486_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__a21o_1 _5566_ (.A1(net13),
    .A2(net61),
    .B1(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__and3_1 _5567_ (.A(net13),
    .B(net61),
    .C(_0500_),
    .X(_0502_));
 sky130_fd_sc_hd__a21oi_1 _5568_ (.A1(_0480_),
    .A2(_0482_),
    .B1(_0483_),
    .Y(_0503_));
 sky130_fd_sc_hd__and3_1 _5569_ (.A(_0480_),
    .B(_0482_),
    .C(_0483_),
    .X(_0504_));
 sky130_fd_sc_hd__or2_1 _5570_ (.A(_0503_),
    .B(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__nand2_1 _5571_ (.A(net10),
    .B(net61),
    .Y(_0507_));
 sky130_fd_sc_hd__xor2_1 _5572_ (.A(_0346_),
    .B(_0348_),
    .X(_0508_));
 sky130_fd_sc_hd__xnor2_1 _5573_ (.A(_0478_),
    .B(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__nand2b_1 _5574_ (.A_N(_0509_),
    .B(_0507_),
    .Y(_0510_));
 sky130_fd_sc_hd__and3_1 _5575_ (.A(net10),
    .B(net61),
    .C(_0509_),
    .X(_0511_));
 sky130_fd_sc_hd__nand2_1 _5576_ (.A(net9),
    .B(net61),
    .Y(_0512_));
 sky130_fd_sc_hd__xor2_1 _5577_ (.A(_0350_),
    .B(_0353_),
    .X(_0513_));
 sky130_fd_sc_hd__xnor2_1 _5578_ (.A(_0477_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__nand2b_1 _5579_ (.A_N(_0514_),
    .B(_0512_),
    .Y(_0515_));
 sky130_fd_sc_hd__and3_1 _5580_ (.A(net9),
    .B(net61),
    .C(_0514_),
    .X(_0516_));
 sky130_fd_sc_hd__nand2_1 _5581_ (.A(net8),
    .B(net61),
    .Y(_0518_));
 sky130_fd_sc_hd__o211ai_2 _5582_ (.A1(_0359_),
    .A2(_0360_),
    .B1(_0367_),
    .C1(_0476_),
    .Y(_0519_));
 sky130_fd_sc_hd__a211o_1 _5583_ (.A1(_0367_),
    .A2(_0476_),
    .B1(_0359_),
    .C1(_0360_),
    .X(_0520_));
 sky130_fd_sc_hd__nand3_1 _5584_ (.A(_0518_),
    .B(_0519_),
    .C(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__a21oi_1 _5585_ (.A1(_0519_),
    .A2(_0520_),
    .B1(_0518_),
    .Y(_0522_));
 sky130_fd_sc_hd__a21o_1 _5586_ (.A1(_0519_),
    .A2(_0520_),
    .B1(_0518_),
    .X(_0523_));
 sky130_fd_sc_hd__and2_1 _5587_ (.A(net7),
    .B(net61),
    .X(_0524_));
 sky130_fd_sc_hd__or2_1 _5588_ (.A(_0366_),
    .B(_0368_),
    .X(_0525_));
 sky130_fd_sc_hd__xnor2_1 _5589_ (.A(_0475_),
    .B(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__and2_1 _5590_ (.A(_0524_),
    .B(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__xor2_1 _5591_ (.A(_0369_),
    .B(_0371_),
    .X(_0529_));
 sky130_fd_sc_hd__nand3_1 _5592_ (.A(_0379_),
    .B(_0474_),
    .C(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__a21o_1 _5593_ (.A1(_0379_),
    .A2(_0474_),
    .B1(_0529_),
    .X(_0531_));
 sky130_fd_sc_hd__and4_1 _5594_ (.A(net6),
    .B(net61),
    .C(_0530_),
    .D(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__a22o_1 _5595_ (.A1(net6),
    .A2(net61),
    .B1(_0530_),
    .B2(_0531_),
    .X(_0533_));
 sky130_fd_sc_hd__nand2_1 _5596_ (.A(net5),
    .B(net61),
    .Y(_0534_));
 sky130_fd_sc_hd__a22o_1 _5597_ (.A1(_0378_),
    .A2(_0379_),
    .B1(_0383_),
    .B2(_0471_),
    .X(_0535_));
 sky130_fd_sc_hd__nand4_1 _5598_ (.A(_0378_),
    .B(_0379_),
    .C(_0383_),
    .D(_0471_),
    .Y(_0536_));
 sky130_fd_sc_hd__a21oi_1 _5599_ (.A1(_0535_),
    .A2(_0536_),
    .B1(_0534_),
    .Y(_0537_));
 sky130_fd_sc_hd__a21o_1 _5600_ (.A1(_0535_),
    .A2(_0536_),
    .B1(_0534_),
    .X(_0538_));
 sky130_fd_sc_hd__and3_1 _5601_ (.A(_0534_),
    .B(_0535_),
    .C(_0536_),
    .X(_0540_));
 sky130_fd_sc_hd__nand2_1 _5602_ (.A(net4),
    .B(net61),
    .Y(_0541_));
 sky130_fd_sc_hd__inv_2 _5603_ (.A(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__xor2_1 _5604_ (.A(_0380_),
    .B(_0382_),
    .X(_0543_));
 sky130_fd_sc_hd__xnor2_2 _5605_ (.A(_0470_),
    .B(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__nor2_1 _5606_ (.A(_0542_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_1 _5607_ (.A(net3),
    .B(net61),
    .Y(_0546_));
 sky130_fd_sc_hd__xor2_1 _5608_ (.A(_0384_),
    .B(_0387_),
    .X(_0547_));
 sky130_fd_sc_hd__xnor2_1 _5609_ (.A(_0469_),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__nand2b_1 _5610_ (.A_N(_0548_),
    .B(_0546_),
    .Y(_0549_));
 sky130_fd_sc_hd__and3_1 _5611_ (.A(net3),
    .B(net61),
    .C(_0548_),
    .X(_0551_));
 sky130_fd_sc_hd__nand2_1 _5612_ (.A(net2),
    .B(net61),
    .Y(_0552_));
 sky130_fd_sc_hd__xor2_1 _5613_ (.A(_0390_),
    .B(_0392_),
    .X(_0553_));
 sky130_fd_sc_hd__nand3_1 _5614_ (.A(_0401_),
    .B(_0468_),
    .C(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__a21o_1 _5615_ (.A1(_0401_),
    .A2(_0468_),
    .B1(_0553_),
    .X(_0555_));
 sky130_fd_sc_hd__a21oi_1 _5616_ (.A1(_0554_),
    .A2(_0555_),
    .B1(_0552_),
    .Y(_0556_));
 sky130_fd_sc_hd__a21o_1 _5617_ (.A1(_0554_),
    .A2(_0555_),
    .B1(_0552_),
    .X(_0557_));
 sky130_fd_sc_hd__and3_1 _5618_ (.A(_0552_),
    .B(_0554_),
    .C(_0555_),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_1 _5619_ (.A(net32),
    .B(net61),
    .Y(_0559_));
 sky130_fd_sc_hd__inv_2 _5620_ (.A(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__and2b_1 _5621_ (.A_N(_0400_),
    .B(_0401_),
    .X(_0562_));
 sky130_fd_sc_hd__xnor2_2 _5622_ (.A(_0467_),
    .B(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__nand2_2 _5623_ (.A(_0560_),
    .B(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2_1 _5624_ (.A(net31),
    .B(net61),
    .Y(_0565_));
 sky130_fd_sc_hd__xor2_1 _5625_ (.A(_0402_),
    .B(_0404_),
    .X(_0566_));
 sky130_fd_sc_hd__xnor2_1 _5626_ (.A(_0466_),
    .B(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__and3_1 _5627_ (.A(net31),
    .B(net61),
    .C(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__nand2b_1 _5628_ (.A_N(_0567_),
    .B(_0565_),
    .Y(_0569_));
 sky130_fd_sc_hd__nand2_1 _5629_ (.A(net30),
    .B(net61),
    .Y(_0570_));
 sky130_fd_sc_hd__xor2_1 _5630_ (.A(_0408_),
    .B(_0410_),
    .X(_0571_));
 sky130_fd_sc_hd__xnor2_1 _5631_ (.A(_0464_),
    .B(_0571_),
    .Y(_0573_));
 sky130_fd_sc_hd__nand2b_1 _5632_ (.A_N(_0573_),
    .B(_0570_),
    .Y(_0574_));
 sky130_fd_sc_hd__and3_1 _5633_ (.A(net30),
    .B(net61),
    .C(_0573_),
    .X(_0575_));
 sky130_fd_sc_hd__nand2_1 _5634_ (.A(net29),
    .B(net61),
    .Y(_0576_));
 sky130_fd_sc_hd__o22ai_1 _5635_ (.A1(_0415_),
    .A2(_0416_),
    .B1(_0422_),
    .B2(_0463_),
    .Y(_0577_));
 sky130_fd_sc_hd__or4_1 _5636_ (.A(_0415_),
    .B(_0416_),
    .C(_0422_),
    .D(_0463_),
    .X(_0578_));
 sky130_fd_sc_hd__a21oi_1 _5637_ (.A1(_0577_),
    .A2(_0578_),
    .B1(_0576_),
    .Y(_0579_));
 sky130_fd_sc_hd__and3_1 _5638_ (.A(_0576_),
    .B(_0577_),
    .C(_0578_),
    .X(_0580_));
 sky130_fd_sc_hd__inv_2 _5639_ (.A(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _5640_ (.A(net28),
    .B(net61),
    .Y(_0582_));
 sky130_fd_sc_hd__inv_2 _5641_ (.A(_0582_),
    .Y(_0584_));
 sky130_fd_sc_hd__xnor2_1 _5642_ (.A(_0419_),
    .B(_0421_),
    .Y(_0585_));
 sky130_fd_sc_hd__xnor2_1 _5643_ (.A(_0461_),
    .B(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__or2_1 _5644_ (.A(_0584_),
    .B(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__nand2_1 _5645_ (.A(net27),
    .B(net61),
    .Y(_0588_));
 sky130_fd_sc_hd__xnor2_1 _5646_ (.A(_0423_),
    .B(_0426_),
    .Y(_0589_));
 sky130_fd_sc_hd__xnor2_1 _5647_ (.A(_0459_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2b_1 _5648_ (.A_N(_0590_),
    .B(_0588_),
    .Y(_0591_));
 sky130_fd_sc_hd__and3_1 _5649_ (.A(net27),
    .B(net61),
    .C(_0590_),
    .X(_0592_));
 sky130_fd_sc_hd__nand2_1 _5650_ (.A(net26),
    .B(net61),
    .Y(_0593_));
 sky130_fd_sc_hd__o21ai_1 _5651_ (.A1(_0431_),
    .A2(_0432_),
    .B1(_0458_),
    .Y(_0595_));
 sky130_fd_sc_hd__or3_1 _5652_ (.A(_0431_),
    .B(_0432_),
    .C(_0458_),
    .X(_0596_));
 sky130_fd_sc_hd__and3_1 _5653_ (.A(_0593_),
    .B(_0595_),
    .C(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__a21oi_1 _5654_ (.A1(_0595_),
    .A2(_0596_),
    .B1(_0593_),
    .Y(_0598_));
 sky130_fd_sc_hd__a2bb2o_1 _5655_ (.A1_N(_0437_),
    .A2_N(_0439_),
    .B1(_0444_),
    .B2(_0457_),
    .X(_0599_));
 sky130_fd_sc_hd__or4bb_1 _5656_ (.A(_0437_),
    .B(_0439_),
    .C_N(_0444_),
    .D_N(_0457_),
    .X(_0600_));
 sky130_fd_sc_hd__nand4_1 _5657_ (.A(net23),
    .B(net61),
    .C(_0599_),
    .D(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__a22oi_1 _5658_ (.A1(net23),
    .A2(net61),
    .B1(_0599_),
    .B2(_0600_),
    .Y(_0602_));
 sky130_fd_sc_hd__a22o_1 _5659_ (.A1(net23),
    .A2(net61),
    .B1(_0599_),
    .B2(_0600_),
    .X(_0603_));
 sky130_fd_sc_hd__nand2_1 _5660_ (.A(net12),
    .B(net61),
    .Y(_0604_));
 sky130_fd_sc_hd__xnor2_1 _5661_ (.A(_0441_),
    .B(_0443_),
    .Y(_0606_));
 sky130_fd_sc_hd__xnor2_2 _5662_ (.A(_0456_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__nand2b_1 _5663_ (.A_N(_0604_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__or2_1 _5664_ (.A(_0448_),
    .B(_0449_),
    .X(_0609_));
 sky130_fd_sc_hd__xnor2_2 _5665_ (.A(_0453_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__nand3_1 _5666_ (.A(net1),
    .B(net61),
    .C(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__o2111ai_4 _5667_ (.A1(net12),
    .A2(_0607_),
    .B1(_0610_),
    .C1(net1),
    .D1(net61),
    .Y(_0612_));
 sky130_fd_sc_hd__a31o_1 _5668_ (.A1(_0601_),
    .A2(_0608_),
    .A3(_0612_),
    .B1(_0602_),
    .X(_0613_));
 sky130_fd_sc_hd__o21bai_2 _5669_ (.A1(_0597_),
    .A2(_0613_),
    .B1_N(_0598_),
    .Y(_0614_));
 sky130_fd_sc_hd__a21o_1 _5670_ (.A1(_0591_),
    .A2(_0614_),
    .B1(_0592_),
    .X(_0615_));
 sky130_fd_sc_hd__a221o_1 _5671_ (.A1(_0584_),
    .A2(_0586_),
    .B1(_0591_),
    .B2(_0614_),
    .C1(_0592_),
    .X(_0617_));
 sky130_fd_sc_hd__a21o_1 _5672_ (.A1(_0587_),
    .A2(_0617_),
    .B1(_0579_),
    .X(_0618_));
 sky130_fd_sc_hd__a31o_2 _5673_ (.A1(_0574_),
    .A2(_0581_),
    .A3(_0618_),
    .B1(_0575_),
    .X(_0619_));
 sky130_fd_sc_hd__o21a_1 _5674_ (.A1(_0568_),
    .A2(_0619_),
    .B1(_0569_),
    .X(_0620_));
 sky130_fd_sc_hd__o221ai_4 _5675_ (.A1(_0560_),
    .A2(_0563_),
    .B1(_0568_),
    .B2(_0619_),
    .C1(_0569_),
    .Y(_0621_));
 sky130_fd_sc_hd__a31oi_4 _5676_ (.A1(_0557_),
    .A2(_0564_),
    .A3(_0621_),
    .B1(_0558_),
    .Y(_0622_));
 sky130_fd_sc_hd__a21oi_1 _5677_ (.A1(_0549_),
    .A2(_0622_),
    .B1(_0551_),
    .Y(_0623_));
 sky130_fd_sc_hd__a221oi_2 _5678_ (.A1(_0542_),
    .A2(_0544_),
    .B1(_0549_),
    .B2(_0622_),
    .C1(_0551_),
    .Y(_0624_));
 sky130_fd_sc_hd__o31ai_2 _5679_ (.A1(_0540_),
    .A2(_0545_),
    .A3(_0624_),
    .B1(_0538_),
    .Y(_0625_));
 sky130_fd_sc_hd__o21a_1 _5680_ (.A1(_0532_),
    .A2(_0625_),
    .B1(_0533_),
    .X(_0626_));
 sky130_fd_sc_hd__o221a_1 _5681_ (.A1(_0524_),
    .A2(_0526_),
    .B1(_0532_),
    .B2(_0625_),
    .C1(_0533_),
    .X(_0628_));
 sky130_fd_sc_hd__o31a_1 _5682_ (.A1(_0522_),
    .A2(_0527_),
    .A3(_0628_),
    .B1(_0521_),
    .X(_0629_));
 sky130_fd_sc_hd__a21o_1 _5683_ (.A1(_0515_),
    .A2(_0629_),
    .B1(_0516_),
    .X(_0630_));
 sky130_fd_sc_hd__a21o_1 _5684_ (.A1(_0510_),
    .A2(_0630_),
    .B1(_0511_),
    .X(_0631_));
 sky130_fd_sc_hd__a2111o_1 _5685_ (.A1(_0510_),
    .A2(_0630_),
    .B1(_0511_),
    .C1(_0503_),
    .D1(_0504_),
    .X(_0632_));
 sky130_fd_sc_hd__and2_1 _5686_ (.A(_0505_),
    .B(_0631_),
    .X(_0633_));
 sky130_fd_sc_hd__nand2_1 _5687_ (.A(net11),
    .B(net61),
    .Y(_0634_));
 sky130_fd_sc_hd__a21bo_1 _5688_ (.A1(_0505_),
    .A2(_0631_),
    .B1_N(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__and3_1 _5689_ (.A(net11),
    .B(net61),
    .C(_0632_),
    .X(_0636_));
 sky130_fd_sc_hd__xor2_1 _5690_ (.A(_0487_),
    .B(_0489_),
    .X(_0637_));
 sky130_fd_sc_hd__xnor2_1 _5691_ (.A(_0492_),
    .B(_0637_),
    .Y(_0639_));
 sky130_fd_sc_hd__a311oi_1 _5692_ (.A1(_0501_),
    .A2(_0632_),
    .A3(_0635_),
    .B1(_0639_),
    .C1(_0502_),
    .Y(_0640_));
 sky130_fd_sc_hd__o311a_1 _5693_ (.A1(_0502_),
    .A2(_0633_),
    .A3(_0636_),
    .B1(_0639_),
    .C1(_0501_),
    .X(_0641_));
 sky130_fd_sc_hd__and2_1 _5694_ (.A(net14),
    .B(net61),
    .X(_0642_));
 sky130_fd_sc_hd__o21ba_1 _5695_ (.A1(_0641_),
    .A2(_0642_),
    .B1_N(_0640_),
    .X(_0643_));
 sky130_fd_sc_hd__o21ai_1 _5696_ (.A1(_0496_),
    .A2(_0643_),
    .B1(_0497_),
    .Y(_0644_));
 sky130_fd_sc_hd__a22oi_2 _5697_ (.A1(net60),
    .A2(_0336_),
    .B1(_0337_),
    .B2(_0493_),
    .Y(_0645_));
 sky130_fd_sc_hd__a21oi_1 _5698_ (.A1(_0644_),
    .A2(_0645_),
    .B1(_3987_),
    .Y(_0646_));
 sky130_fd_sc_hd__a21oi_1 _5699_ (.A1(net62),
    .A2(_1716_),
    .B1(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2_1 _5700_ (.A(net62),
    .B(_0646_),
    .Y(_0648_));
 sky130_fd_sc_hd__and2b_1 _5701_ (.A_N(_0647_),
    .B(_0648_),
    .X(_0650_));
 sky130_fd_sc_hd__xor2_1 _5702_ (.A(_0644_),
    .B(_0645_),
    .X(_0651_));
 sky130_fd_sc_hd__xnor2_1 _5703_ (.A(_3987_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__nand2_1 _5704_ (.A(net14),
    .B(net62),
    .Y(_0653_));
 sky130_fd_sc_hd__xor2_1 _5705_ (.A(_3988_),
    .B(_0494_),
    .X(_0654_));
 sky130_fd_sc_hd__xnor2_1 _5706_ (.A(_0643_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__nand2b_1 _5707_ (.A_N(_0655_),
    .B(_0653_),
    .Y(_0656_));
 sky130_fd_sc_hd__and3_1 _5708_ (.A(net14),
    .B(net62),
    .C(_0655_),
    .X(_0657_));
 sky130_fd_sc_hd__nand2_1 _5709_ (.A(net11),
    .B(net62),
    .Y(_0658_));
 sky130_fd_sc_hd__xor2_1 _5710_ (.A(_0498_),
    .B(_0500_),
    .X(_0659_));
 sky130_fd_sc_hd__o21ai_1 _5711_ (.A1(_0633_),
    .A2(_0636_),
    .B1(_0659_),
    .Y(_0661_));
 sky130_fd_sc_hd__or3_1 _5712_ (.A(_0633_),
    .B(_0636_),
    .C(_0659_),
    .X(_0662_));
 sky130_fd_sc_hd__a21oi_1 _5713_ (.A1(_0661_),
    .A2(_0662_),
    .B1(_0658_),
    .Y(_0663_));
 sky130_fd_sc_hd__and3_1 _5714_ (.A(_0658_),
    .B(_0661_),
    .C(_0662_),
    .X(_0664_));
 sky130_fd_sc_hd__nand3_1 _5715_ (.A(_0658_),
    .B(_0661_),
    .C(_0662_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand2_1 _5716_ (.A(net9),
    .B(net62),
    .Y(_0666_));
 sky130_fd_sc_hd__xor2_1 _5717_ (.A(_0507_),
    .B(_0509_),
    .X(_0667_));
 sky130_fd_sc_hd__xnor2_1 _5718_ (.A(_0630_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__and3_1 _5719_ (.A(net9),
    .B(net62),
    .C(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__nand2b_1 _5720_ (.A_N(_0668_),
    .B(_0666_),
    .Y(_0670_));
 sky130_fd_sc_hd__nand2_1 _5721_ (.A(net8),
    .B(net62),
    .Y(_0672_));
 sky130_fd_sc_hd__xor2_1 _5722_ (.A(_0512_),
    .B(_0514_),
    .X(_0673_));
 sky130_fd_sc_hd__xnor2_1 _5723_ (.A(_0629_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__a21o_1 _5724_ (.A1(net8),
    .A2(net62),
    .B1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__and3_1 _5725_ (.A(net8),
    .B(net62),
    .C(_0674_),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_1 _5726_ (.A(net7),
    .B(net62),
    .Y(_0677_));
 sky130_fd_sc_hd__inv_2 _5727_ (.A(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__o211ai_2 _5728_ (.A1(_0527_),
    .A2(_0628_),
    .B1(_0521_),
    .C1(_0523_),
    .Y(_0679_));
 sky130_fd_sc_hd__a211o_1 _5729_ (.A1(_0521_),
    .A2(_0523_),
    .B1(_0527_),
    .C1(_0628_),
    .X(_0680_));
 sky130_fd_sc_hd__a21oi_1 _5730_ (.A1(_0679_),
    .A2(_0680_),
    .B1(_0678_),
    .Y(_0681_));
 sky130_fd_sc_hd__a21o_1 _5731_ (.A1(_0679_),
    .A2(_0680_),
    .B1(_0678_),
    .X(_0683_));
 sky130_fd_sc_hd__and3_1 _5732_ (.A(_0678_),
    .B(_0679_),
    .C(_0680_),
    .X(_0684_));
 sky130_fd_sc_hd__nand2_1 _5733_ (.A(net6),
    .B(net62),
    .Y(_0685_));
 sky130_fd_sc_hd__xnor2_1 _5734_ (.A(_0524_),
    .B(_0526_),
    .Y(_0686_));
 sky130_fd_sc_hd__xnor2_1 _5735_ (.A(_0626_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__and3_1 _5736_ (.A(net6),
    .B(net62),
    .C(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__a21o_1 _5737_ (.A1(net6),
    .A2(net62),
    .B1(_0687_),
    .X(_0689_));
 sky130_fd_sc_hd__and2_1 _5738_ (.A(net5),
    .B(net62),
    .X(_0690_));
 sky130_fd_sc_hd__nand2b_1 _5739_ (.A_N(_0532_),
    .B(_0533_),
    .Y(_0691_));
 sky130_fd_sc_hd__xnor2_1 _5740_ (.A(_0625_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__or2_1 _5741_ (.A(_0690_),
    .B(_0692_),
    .X(_0694_));
 sky130_fd_sc_hd__nand2_1 _5742_ (.A(net4),
    .B(net62),
    .Y(_0695_));
 sky130_fd_sc_hd__o22a_1 _5743_ (.A1(_0537_),
    .A2(_0540_),
    .B1(_0545_),
    .B2(_0624_),
    .X(_0696_));
 sky130_fd_sc_hd__or4_1 _5744_ (.A(_0537_),
    .B(_0540_),
    .C(_0545_),
    .D(_0624_),
    .X(_0697_));
 sky130_fd_sc_hd__and2b_1 _5745_ (.A_N(_0696_),
    .B(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__and3_1 _5746_ (.A(net4),
    .B(net62),
    .C(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__a21o_1 _5747_ (.A1(net4),
    .A2(net62),
    .B1(_0698_),
    .X(_0700_));
 sky130_fd_sc_hd__nand2_1 _5748_ (.A(net3),
    .B(net62),
    .Y(_0701_));
 sky130_fd_sc_hd__xnor2_1 _5749_ (.A(_0541_),
    .B(_0544_),
    .Y(_0702_));
 sky130_fd_sc_hd__xnor2_2 _5750_ (.A(_0623_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__a21oi_1 _5751_ (.A1(net3),
    .A2(net62),
    .B1(_0703_),
    .Y(_0705_));
 sky130_fd_sc_hd__nand2b_1 _5752_ (.A_N(_0701_),
    .B(_0703_),
    .Y(_0706_));
 sky130_fd_sc_hd__nand2_1 _5753_ (.A(net2),
    .B(net62),
    .Y(_0707_));
 sky130_fd_sc_hd__xor2_1 _5754_ (.A(_0546_),
    .B(_0548_),
    .X(_0708_));
 sky130_fd_sc_hd__xnor2_2 _5755_ (.A(_0622_),
    .B(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__and2b_1 _5756_ (.A_N(_0709_),
    .B(_0707_),
    .X(_0710_));
 sky130_fd_sc_hd__nand2b_1 _5757_ (.A_N(_0707_),
    .B(_0709_),
    .Y(_0711_));
 sky130_fd_sc_hd__o211ai_2 _5758_ (.A1(_0556_),
    .A2(_0558_),
    .B1(_0564_),
    .C1(_0621_),
    .Y(_0712_));
 sky130_fd_sc_hd__a211o_1 _5759_ (.A1(_0564_),
    .A2(_0621_),
    .B1(_0556_),
    .C1(_0558_),
    .X(_0713_));
 sky130_fd_sc_hd__and2_1 _5760_ (.A(net32),
    .B(net62),
    .X(_0714_));
 sky130_fd_sc_hd__a21oi_1 _5761_ (.A1(_0712_),
    .A2(_0713_),
    .B1(_0714_),
    .Y(_0716_));
 sky130_fd_sc_hd__and3_1 _5762_ (.A(_0712_),
    .B(_0713_),
    .C(_0714_),
    .X(_0717_));
 sky130_fd_sc_hd__nand3_1 _5763_ (.A(_0712_),
    .B(_0713_),
    .C(_0714_),
    .Y(_0718_));
 sky130_fd_sc_hd__nand2_1 _5764_ (.A(net31),
    .B(net62),
    .Y(_0719_));
 sky130_fd_sc_hd__xnor2_1 _5765_ (.A(_0559_),
    .B(_0563_),
    .Y(_0720_));
 sky130_fd_sc_hd__xnor2_1 _5766_ (.A(_0620_),
    .B(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__or2_1 _5767_ (.A(_0719_),
    .B(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__nand2_1 _5768_ (.A(net30),
    .B(net62),
    .Y(_0723_));
 sky130_fd_sc_hd__xor2_1 _5769_ (.A(_0565_),
    .B(_0567_),
    .X(_0724_));
 sky130_fd_sc_hd__xnor2_2 _5770_ (.A(_0619_),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__nand2b_1 _5771_ (.A_N(_0723_),
    .B(_0725_),
    .Y(_0727_));
 sky130_fd_sc_hd__a21oi_1 _5772_ (.A1(net30),
    .A2(net62),
    .B1(_0725_),
    .Y(_0728_));
 sky130_fd_sc_hd__xor2_1 _5773_ (.A(_0570_),
    .B(_0573_),
    .X(_0729_));
 sky130_fd_sc_hd__a21bo_1 _5774_ (.A1(_0581_),
    .A2(_0618_),
    .B1_N(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__or3b_1 _5775_ (.A(_0580_),
    .B(_0729_),
    .C_N(_0618_),
    .X(_0731_));
 sky130_fd_sc_hd__a22oi_1 _5776_ (.A1(net29),
    .A2(net62),
    .B1(_0730_),
    .B2(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__a22o_1 _5777_ (.A1(net29),
    .A2(net62),
    .B1(_0730_),
    .B2(_0731_),
    .X(_0733_));
 sky130_fd_sc_hd__and4_1 _5778_ (.A(net29),
    .B(net62),
    .C(_0730_),
    .D(_0731_),
    .X(_0734_));
 sky130_fd_sc_hd__nand2_1 _5779_ (.A(net28),
    .B(net62),
    .Y(_0735_));
 sky130_fd_sc_hd__o211ai_2 _5780_ (.A1(_0579_),
    .A2(_0580_),
    .B1(_0587_),
    .C1(_0617_),
    .Y(_0736_));
 sky130_fd_sc_hd__a211o_1 _5781_ (.A1(_0587_),
    .A2(_0617_),
    .B1(_0579_),
    .C1(_0580_),
    .X(_0738_));
 sky130_fd_sc_hd__a21oi_1 _5782_ (.A1(_0736_),
    .A2(_0738_),
    .B1(_0735_),
    .Y(_0739_));
 sky130_fd_sc_hd__a21o_1 _5783_ (.A1(_0736_),
    .A2(_0738_),
    .B1(_0735_),
    .X(_0740_));
 sky130_fd_sc_hd__and3_1 _5784_ (.A(_0735_),
    .B(_0736_),
    .C(_0738_),
    .X(_0741_));
 sky130_fd_sc_hd__nand2_1 _5785_ (.A(net27),
    .B(net62),
    .Y(_0742_));
 sky130_fd_sc_hd__xnor2_1 _5786_ (.A(_0582_),
    .B(_0586_),
    .Y(_0743_));
 sky130_fd_sc_hd__xnor2_1 _5787_ (.A(_0615_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__or2_1 _5788_ (.A(_0742_),
    .B(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__nand2_1 _5789_ (.A(net26),
    .B(net62),
    .Y(_0746_));
 sky130_fd_sc_hd__xor2_1 _5790_ (.A(_0588_),
    .B(_0590_),
    .X(_0747_));
 sky130_fd_sc_hd__xnor2_1 _5791_ (.A(_0614_),
    .B(_0747_),
    .Y(_0749_));
 sky130_fd_sc_hd__a21oi_1 _5792_ (.A1(net26),
    .A2(net62),
    .B1(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__nand2b_1 _5793_ (.A_N(_0746_),
    .B(_0749_),
    .Y(_0751_));
 sky130_fd_sc_hd__o21ai_1 _5794_ (.A1(_0597_),
    .A2(_0598_),
    .B1(_0613_),
    .Y(_0752_));
 sky130_fd_sc_hd__or3_1 _5795_ (.A(_0597_),
    .B(_0598_),
    .C(_0613_),
    .X(_0753_));
 sky130_fd_sc_hd__and4_1 _5796_ (.A(net23),
    .B(net62),
    .C(_0752_),
    .D(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__a22oi_2 _5797_ (.A1(net23),
    .A2(net62),
    .B1(_0752_),
    .B2(_0753_),
    .Y(_0755_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(net12),
    .B(net62),
    .Y(_0756_));
 sky130_fd_sc_hd__nand4_1 _5799_ (.A(_0601_),
    .B(_0603_),
    .C(_0608_),
    .D(_0612_),
    .Y(_0757_));
 sky130_fd_sc_hd__a22o_1 _5800_ (.A1(_0601_),
    .A2(_0603_),
    .B1(_0608_),
    .B2(_0612_),
    .X(_0758_));
 sky130_fd_sc_hd__a21oi_1 _5801_ (.A1(_0757_),
    .A2(_0758_),
    .B1(_0756_),
    .Y(_0760_));
 sky130_fd_sc_hd__a21o_1 _5802_ (.A1(_0757_),
    .A2(_0758_),
    .B1(_0756_),
    .X(_0761_));
 sky130_fd_sc_hd__and3_1 _5803_ (.A(_0756_),
    .B(_0757_),
    .C(_0758_),
    .X(_0762_));
 sky130_fd_sc_hd__xor2_1 _5804_ (.A(_0604_),
    .B(_0607_),
    .X(_0763_));
 sky130_fd_sc_hd__a21oi_1 _5805_ (.A1(_0611_),
    .A2(_0763_),
    .B1(_4198_),
    .Y(_0764_));
 sky130_fd_sc_hd__o211ai_2 _5806_ (.A1(_0611_),
    .A2(_0763_),
    .B1(_0764_),
    .C1(net62),
    .Y(_0765_));
 sky130_fd_sc_hd__a21o_1 _5807_ (.A1(_0761_),
    .A2(_0765_),
    .B1(_0762_),
    .X(_0766_));
 sky130_fd_sc_hd__a21oi_1 _5808_ (.A1(_0761_),
    .A2(_0765_),
    .B1(_0762_),
    .Y(_0767_));
 sky130_fd_sc_hd__o21bai_2 _5809_ (.A1(_0754_),
    .A2(_0767_),
    .B1_N(_0755_),
    .Y(_0768_));
 sky130_fd_sc_hd__a21oi_1 _5810_ (.A1(_0751_),
    .A2(_0768_),
    .B1(_0750_),
    .Y(_0769_));
 sky130_fd_sc_hd__a221o_1 _5811_ (.A1(_0742_),
    .A2(_0744_),
    .B1(_0751_),
    .B2(_0768_),
    .C1(_0750_),
    .X(_0771_));
 sky130_fd_sc_hd__a31oi_1 _5812_ (.A1(_0740_),
    .A2(_0745_),
    .A3(_0771_),
    .B1(_0741_),
    .Y(_0772_));
 sky130_fd_sc_hd__a21oi_1 _5813_ (.A1(_0733_),
    .A2(_0772_),
    .B1(_0734_),
    .Y(_0773_));
 sky130_fd_sc_hd__a21oi_1 _5814_ (.A1(_0727_),
    .A2(_0773_),
    .B1(_0728_),
    .Y(_0774_));
 sky130_fd_sc_hd__a221o_1 _5815_ (.A1(_0719_),
    .A2(_0721_),
    .B1(_0727_),
    .B2(_0773_),
    .C1(_0728_),
    .X(_0775_));
 sky130_fd_sc_hd__a21o_1 _5816_ (.A1(_0722_),
    .A2(_0775_),
    .B1(_0716_),
    .X(_0776_));
 sky130_fd_sc_hd__a31o_1 _5817_ (.A1(_0711_),
    .A2(_0718_),
    .A3(_0776_),
    .B1(_0710_),
    .X(_0777_));
 sky130_fd_sc_hd__o21ai_2 _5818_ (.A1(_0705_),
    .A2(_0777_),
    .B1(_0706_),
    .Y(_0778_));
 sky130_fd_sc_hd__a21o_1 _5819_ (.A1(_0700_),
    .A2(_0778_),
    .B1(_0699_),
    .X(_0779_));
 sky130_fd_sc_hd__a221o_1 _5820_ (.A1(_0690_),
    .A2(_0692_),
    .B1(_0700_),
    .B2(_0778_),
    .C1(_0699_),
    .X(_0780_));
 sky130_fd_sc_hd__a31o_1 _5821_ (.A1(_0689_),
    .A2(_0694_),
    .A3(_0780_),
    .B1(_0688_),
    .X(_0782_));
 sky130_fd_sc_hd__a311o_1 _5822_ (.A1(_0689_),
    .A2(_0694_),
    .A3(_0780_),
    .B1(_0688_),
    .C1(_0684_),
    .X(_0783_));
 sky130_fd_sc_hd__a31o_1 _5823_ (.A1(_0675_),
    .A2(_0683_),
    .A3(_0783_),
    .B1(_0676_),
    .X(_0784_));
 sky130_fd_sc_hd__o21a_1 _5824_ (.A1(_0669_),
    .A2(_0784_),
    .B1(_0670_),
    .X(_0785_));
 sky130_fd_sc_hd__xor2_1 _5825_ (.A(_0505_),
    .B(_0631_),
    .X(_0786_));
 sky130_fd_sc_hd__xnor2_1 _5826_ (.A(_0634_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__or2_1 _5827_ (.A(_0785_),
    .B(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_1 _5828_ (.A(net10),
    .B(net62),
    .Y(_0789_));
 sky130_fd_sc_hd__a21bo_1 _5829_ (.A1(_0785_),
    .A2(_0787_),
    .B1_N(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__a31o_1 _5830_ (.A1(_0665_),
    .A2(_0788_),
    .A3(_0790_),
    .B1(_0663_),
    .X(_0791_));
 sky130_fd_sc_hd__nor2_1 _5831_ (.A(_0640_),
    .B(_0641_),
    .Y(_0793_));
 sky130_fd_sc_hd__xor2_1 _5832_ (.A(_0642_),
    .B(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__or2_1 _5833_ (.A(_0791_),
    .B(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__nand2_1 _5834_ (.A(net13),
    .B(net62),
    .Y(_0796_));
 sky130_fd_sc_hd__a21bo_1 _5835_ (.A1(_0791_),
    .A2(_0794_),
    .B1_N(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__a31o_1 _5836_ (.A1(_0656_),
    .A2(_0795_),
    .A3(_0797_),
    .B1(_0657_),
    .X(_0798_));
 sky130_fd_sc_hd__nand2_1 _5837_ (.A(_0652_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__nand2_1 _5838_ (.A(net15),
    .B(net62),
    .Y(_0800_));
 sky130_fd_sc_hd__o21bai_1 _5839_ (.A1(_0652_),
    .A2(_0798_),
    .B1_N(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__a21o_1 _5840_ (.A1(_0799_),
    .A2(_0801_),
    .B1(_0650_),
    .X(_0802_));
 sky130_fd_sc_hd__nand3_1 _5841_ (.A(_0650_),
    .B(_0799_),
    .C(_0801_),
    .Y(_0804_));
 sky130_fd_sc_hd__a21oi_1 _5842_ (.A1(_0802_),
    .A2(_0804_),
    .B1(_3986_),
    .Y(_0805_));
 sky130_fd_sc_hd__a21o_1 _5843_ (.A1(_0802_),
    .A2(_0804_),
    .B1(_3986_),
    .X(_0806_));
 sky130_fd_sc_hd__nand3_1 _5844_ (.A(_3986_),
    .B(_0802_),
    .C(_0804_),
    .Y(_0807_));
 sky130_fd_sc_hd__xnor2_1 _5845_ (.A(_0653_),
    .B(_0655_),
    .Y(_0808_));
 sky130_fd_sc_hd__a21o_1 _5846_ (.A1(_0795_),
    .A2(_0797_),
    .B1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__nand3_1 _5847_ (.A(_0795_),
    .B(_0797_),
    .C(_0808_),
    .Y(_0810_));
 sky130_fd_sc_hd__a22o_1 _5848_ (.A1(net13),
    .A2(net63),
    .B1(_0809_),
    .B2(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__and4_1 _5849_ (.A(net13),
    .B(net63),
    .C(_0809_),
    .D(_0810_),
    .X(_0812_));
 sky130_fd_sc_hd__nand4_1 _5850_ (.A(net13),
    .B(net63),
    .C(_0809_),
    .D(_0810_),
    .Y(_0813_));
 sky130_fd_sc_hd__and2_1 _5851_ (.A(net10),
    .B(net63),
    .X(_0815_));
 sky130_fd_sc_hd__a2bb2o_1 _5852_ (.A1_N(_0663_),
    .A2_N(_0664_),
    .B1(_0788_),
    .B2(_0790_),
    .X(_0816_));
 sky130_fd_sc_hd__or4bb_1 _5853_ (.A(_0663_),
    .B(_0664_),
    .C_N(_0788_),
    .D_N(_0790_),
    .X(_0817_));
 sky130_fd_sc_hd__a21oi_1 _5854_ (.A1(_0816_),
    .A2(_0817_),
    .B1(_0815_),
    .Y(_0818_));
 sky130_fd_sc_hd__a21o_1 _5855_ (.A1(_0816_),
    .A2(_0817_),
    .B1(_0815_),
    .X(_0819_));
 sky130_fd_sc_hd__and3_1 _5856_ (.A(_0815_),
    .B(_0816_),
    .C(_0817_),
    .X(_0820_));
 sky130_fd_sc_hd__nand2_1 _5857_ (.A(net8),
    .B(net63),
    .Y(_0821_));
 sky130_fd_sc_hd__xor2_1 _5858_ (.A(_0666_),
    .B(_0668_),
    .X(_0822_));
 sky130_fd_sc_hd__xnor2_1 _5859_ (.A(_0784_),
    .B(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__a21o_1 _5860_ (.A1(net8),
    .A2(net63),
    .B1(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__and3_1 _5861_ (.A(net8),
    .B(net63),
    .C(_0823_),
    .X(_0826_));
 sky130_fd_sc_hd__and2_1 _5862_ (.A(net7),
    .B(net63),
    .X(_0827_));
 sky130_fd_sc_hd__xnor2_1 _5863_ (.A(_0672_),
    .B(_0674_),
    .Y(_0828_));
 sky130_fd_sc_hd__a21o_1 _5864_ (.A1(_0683_),
    .A2(_0783_),
    .B1(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__nand3_1 _5865_ (.A(_0683_),
    .B(_0783_),
    .C(_0828_),
    .Y(_0830_));
 sky130_fd_sc_hd__nand2_1 _5866_ (.A(_0829_),
    .B(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__a21o_1 _5867_ (.A1(_0829_),
    .A2(_0830_),
    .B1(_0827_),
    .X(_0832_));
 sky130_fd_sc_hd__and3_1 _5868_ (.A(_0827_),
    .B(_0829_),
    .C(_0830_),
    .X(_0833_));
 sky130_fd_sc_hd__nand2_1 _5869_ (.A(net6),
    .B(net63),
    .Y(_0834_));
 sky130_fd_sc_hd__or2_1 _5870_ (.A(_0681_),
    .B(_0684_),
    .X(_0835_));
 sky130_fd_sc_hd__xnor2_1 _5871_ (.A(_0782_),
    .B(_0835_),
    .Y(_0837_));
 sky130_fd_sc_hd__nand2b_1 _5872_ (.A_N(_0837_),
    .B(_0834_),
    .Y(_0838_));
 sky130_fd_sc_hd__and3_1 _5873_ (.A(net6),
    .B(net63),
    .C(_0837_),
    .X(_0839_));
 sky130_fd_sc_hd__and2_1 _5874_ (.A(net5),
    .B(net63),
    .X(_0840_));
 sky130_fd_sc_hd__xnor2_1 _5875_ (.A(_0685_),
    .B(_0687_),
    .Y(_0841_));
 sky130_fd_sc_hd__a21o_1 _5876_ (.A1(_0694_),
    .A2(_0780_),
    .B1(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__nand3_1 _5877_ (.A(_0694_),
    .B(_0780_),
    .C(_0841_),
    .Y(_0843_));
 sky130_fd_sc_hd__a21o_1 _5878_ (.A1(_0842_),
    .A2(_0843_),
    .B1(_0840_),
    .X(_0844_));
 sky130_fd_sc_hd__and3_1 _5879_ (.A(_0840_),
    .B(_0842_),
    .C(_0843_),
    .X(_0845_));
 sky130_fd_sc_hd__nand3_1 _5880_ (.A(_0840_),
    .B(_0842_),
    .C(_0843_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _5881_ (.A(net4),
    .B(net63),
    .Y(_0848_));
 sky130_fd_sc_hd__inv_2 _5882_ (.A(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__xnor2_1 _5883_ (.A(_0690_),
    .B(_0692_),
    .Y(_0850_));
 sky130_fd_sc_hd__xnor2_1 _5884_ (.A(_0779_),
    .B(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__or2_1 _5885_ (.A(_0849_),
    .B(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__nand2_1 _5886_ (.A(net3),
    .B(net63),
    .Y(_0853_));
 sky130_fd_sc_hd__xor2_1 _5887_ (.A(_0695_),
    .B(_0698_),
    .X(_0854_));
 sky130_fd_sc_hd__xnor2_1 _5888_ (.A(_0778_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__and3_1 _5889_ (.A(net3),
    .B(net63),
    .C(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__a21o_1 _5890_ (.A1(net3),
    .A2(net63),
    .B1(_0855_),
    .X(_0857_));
 sky130_fd_sc_hd__nand2_1 _5891_ (.A(net2),
    .B(net63),
    .Y(_0859_));
 sky130_fd_sc_hd__xnor2_1 _5892_ (.A(_0701_),
    .B(_0703_),
    .Y(_0860_));
 sky130_fd_sc_hd__xnor2_1 _5893_ (.A(_0777_),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__nand2b_1 _5894_ (.A_N(_0861_),
    .B(_0859_),
    .Y(_0862_));
 sky130_fd_sc_hd__and3_1 _5895_ (.A(net2),
    .B(net63),
    .C(_0861_),
    .X(_0863_));
 sky130_fd_sc_hd__xor2_1 _5896_ (.A(_0707_),
    .B(_0709_),
    .X(_0864_));
 sky130_fd_sc_hd__a21o_1 _5897_ (.A1(_0718_),
    .A2(_0776_),
    .B1(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__nand3_1 _5898_ (.A(_0718_),
    .B(_0776_),
    .C(_0864_),
    .Y(_0866_));
 sky130_fd_sc_hd__a22o_1 _5899_ (.A1(net32),
    .A2(net63),
    .B1(_0865_),
    .B2(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__and4_1 _5900_ (.A(net32),
    .B(net63),
    .C(_0865_),
    .D(_0866_),
    .X(_0868_));
 sky130_fd_sc_hd__nand4_1 _5901_ (.A(net32),
    .B(net63),
    .C(_0865_),
    .D(_0866_),
    .Y(_0870_));
 sky130_fd_sc_hd__o211ai_2 _5902_ (.A1(_0716_),
    .A2(_0717_),
    .B1(_0722_),
    .C1(_0775_),
    .Y(_0871_));
 sky130_fd_sc_hd__a211o_1 _5903_ (.A1(_0722_),
    .A2(_0775_),
    .B1(_0716_),
    .C1(_0717_),
    .X(_0872_));
 sky130_fd_sc_hd__and4_1 _5904_ (.A(net31),
    .B(net63),
    .C(_0871_),
    .D(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__a22oi_1 _5905_ (.A1(net31),
    .A2(net63),
    .B1(_0871_),
    .B2(_0872_),
    .Y(_0874_));
 sky130_fd_sc_hd__a22o_1 _5906_ (.A1(net31),
    .A2(net63),
    .B1(_0871_),
    .B2(_0872_),
    .X(_0875_));
 sky130_fd_sc_hd__nand2_1 _5907_ (.A(net30),
    .B(net63),
    .Y(_0876_));
 sky130_fd_sc_hd__inv_2 _5908_ (.A(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__xnor2_1 _5909_ (.A(_0719_),
    .B(_0721_),
    .Y(_0878_));
 sky130_fd_sc_hd__xnor2_1 _5910_ (.A(_0774_),
    .B(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__or2_1 _5911_ (.A(_0877_),
    .B(_0879_),
    .X(_0881_));
 sky130_fd_sc_hd__nand2_1 _5912_ (.A(net29),
    .B(net63),
    .Y(_0882_));
 sky130_fd_sc_hd__xnor2_1 _5913_ (.A(_0723_),
    .B(_0725_),
    .Y(_0883_));
 sky130_fd_sc_hd__xnor2_1 _5914_ (.A(_0773_),
    .B(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__a21o_1 _5915_ (.A1(net29),
    .A2(net63),
    .B1(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__and3_1 _5916_ (.A(net29),
    .B(net63),
    .C(_0884_),
    .X(_0886_));
 sky130_fd_sc_hd__nand2_1 _5917_ (.A(net28),
    .B(net63),
    .Y(_0887_));
 sky130_fd_sc_hd__o21ai_1 _5918_ (.A1(_0732_),
    .A2(_0734_),
    .B1(_0772_),
    .Y(_0888_));
 sky130_fd_sc_hd__or3b_1 _5919_ (.A(_0772_),
    .B(_0734_),
    .C_N(_0733_),
    .X(_0889_));
 sky130_fd_sc_hd__nand3_1 _5920_ (.A(_0887_),
    .B(_0888_),
    .C(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__a21o_1 _5921_ (.A1(_0888_),
    .A2(_0889_),
    .B1(_0887_),
    .X(_0892_));
 sky130_fd_sc_hd__and2_1 _5922_ (.A(net27),
    .B(net63),
    .X(_0893_));
 sky130_fd_sc_hd__o211ai_2 _5923_ (.A1(_0739_),
    .A2(_0741_),
    .B1(_0745_),
    .C1(_0771_),
    .Y(_0894_));
 sky130_fd_sc_hd__a211o_1 _5924_ (.A1(_0745_),
    .A2(_0771_),
    .B1(_0739_),
    .C1(_0741_),
    .X(_0895_));
 sky130_fd_sc_hd__and3_1 _5925_ (.A(_0893_),
    .B(_0894_),
    .C(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__a21oi_1 _5926_ (.A1(_0894_),
    .A2(_0895_),
    .B1(_0893_),
    .Y(_0897_));
 sky130_fd_sc_hd__a21o_1 _5927_ (.A1(_0894_),
    .A2(_0895_),
    .B1(_0893_),
    .X(_0898_));
 sky130_fd_sc_hd__nand2_1 _5928_ (.A(net26),
    .B(net63),
    .Y(_0899_));
 sky130_fd_sc_hd__inv_2 _5929_ (.A(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__xnor2_1 _5930_ (.A(_0742_),
    .B(_0744_),
    .Y(_0901_));
 sky130_fd_sc_hd__xnor2_1 _5931_ (.A(_0769_),
    .B(_0901_),
    .Y(_0903_));
 sky130_fd_sc_hd__and2_1 _5932_ (.A(_0900_),
    .B(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__nand2_1 _5933_ (.A(net23),
    .B(net63),
    .Y(_0905_));
 sky130_fd_sc_hd__xnor2_1 _5934_ (.A(_0746_),
    .B(_0749_),
    .Y(_0906_));
 sky130_fd_sc_hd__xnor2_1 _5935_ (.A(_0768_),
    .B(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__and3_1 _5936_ (.A(net23),
    .B(net63),
    .C(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__a21o_1 _5937_ (.A1(net23),
    .A2(net63),
    .B1(_0907_),
    .X(_0909_));
 sky130_fd_sc_hd__o21ai_1 _5938_ (.A1(_0754_),
    .A2(_0755_),
    .B1(_0766_),
    .Y(_0910_));
 sky130_fd_sc_hd__or3_1 _5939_ (.A(_0754_),
    .B(_0755_),
    .C(_0766_),
    .X(_0911_));
 sky130_fd_sc_hd__a22o_1 _5940_ (.A1(net12),
    .A2(net63),
    .B1(_0910_),
    .B2(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__nand4_2 _5941_ (.A(net12),
    .B(net63),
    .C(_0910_),
    .D(_0911_),
    .Y(_0914_));
 sky130_fd_sc_hd__nor2_1 _5942_ (.A(_0760_),
    .B(_0762_),
    .Y(_0915_));
 sky130_fd_sc_hd__xor2_1 _5943_ (.A(_0765_),
    .B(_0915_),
    .X(_0916_));
 sky130_fd_sc_hd__or3b_1 _5944_ (.A(_4198_),
    .B(_0916_),
    .C_N(net63),
    .X(_0917_));
 sky130_fd_sc_hd__a21boi_2 _5945_ (.A1(_0914_),
    .A2(_0917_),
    .B1_N(_0912_),
    .Y(_0918_));
 sky130_fd_sc_hd__o21ai_1 _5946_ (.A1(_0908_),
    .A2(_0918_),
    .B1(_0909_),
    .Y(_0919_));
 sky130_fd_sc_hd__o221a_1 _5947_ (.A1(_0900_),
    .A2(_0903_),
    .B1(_0908_),
    .B2(_0918_),
    .C1(_0909_),
    .X(_0920_));
 sky130_fd_sc_hd__o31a_1 _5948_ (.A1(_0896_),
    .A2(_0904_),
    .A3(_0920_),
    .B1(_0898_),
    .X(_0921_));
 sky130_fd_sc_hd__a21bo_1 _5949_ (.A1(_0890_),
    .A2(_0921_),
    .B1_N(_0892_),
    .X(_0922_));
 sky130_fd_sc_hd__a21oi_1 _5950_ (.A1(_0885_),
    .A2(_0922_),
    .B1(_0886_),
    .Y(_0923_));
 sky130_fd_sc_hd__a221o_1 _5951_ (.A1(_0877_),
    .A2(_0879_),
    .B1(_0885_),
    .B2(_0922_),
    .C1(_0886_),
    .X(_0925_));
 sky130_fd_sc_hd__a21o_1 _5952_ (.A1(_0881_),
    .A2(_0925_),
    .B1(_0873_),
    .X(_0926_));
 sky130_fd_sc_hd__a31o_1 _5953_ (.A1(_0867_),
    .A2(_0875_),
    .A3(_0926_),
    .B1(_0868_),
    .X(_0927_));
 sky130_fd_sc_hd__a21o_1 _5954_ (.A1(_0862_),
    .A2(_0927_),
    .B1(_0863_),
    .X(_0928_));
 sky130_fd_sc_hd__a21oi_1 _5955_ (.A1(_0857_),
    .A2(_0928_),
    .B1(_0856_),
    .Y(_0929_));
 sky130_fd_sc_hd__a221o_1 _5956_ (.A1(_0849_),
    .A2(_0851_),
    .B1(_0857_),
    .B2(_0928_),
    .C1(_0856_),
    .X(_0930_));
 sky130_fd_sc_hd__and3_1 _5957_ (.A(_0844_),
    .B(_0852_),
    .C(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__a31o_1 _5958_ (.A1(_0844_),
    .A2(_0852_),
    .A3(_0930_),
    .B1(_0845_),
    .X(_0932_));
 sky130_fd_sc_hd__a21o_1 _5959_ (.A1(_0838_),
    .A2(_0932_),
    .B1(_0839_),
    .X(_0933_));
 sky130_fd_sc_hd__o311a_1 _5960_ (.A1(_0839_),
    .A2(_0845_),
    .A3(_0931_),
    .B1(_0838_),
    .C1(_0832_),
    .X(_0934_));
 sky130_fd_sc_hd__o31a_1 _5961_ (.A1(_0826_),
    .A2(_0833_),
    .A3(_0934_),
    .B1(_0824_),
    .X(_0936_));
 sky130_fd_sc_hd__xor2_1 _5962_ (.A(_0785_),
    .B(_0787_),
    .X(_0937_));
 sky130_fd_sc_hd__xnor2_1 _5963_ (.A(_0789_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__or2_1 _5964_ (.A(_0936_),
    .B(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__nand2_1 _5965_ (.A(net9),
    .B(net63),
    .Y(_0940_));
 sky130_fd_sc_hd__a21bo_1 _5966_ (.A1(_0936_),
    .A2(_0938_),
    .B1_N(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__a31o_1 _5967_ (.A1(_0819_),
    .A2(_0939_),
    .A3(_0941_),
    .B1(_0820_),
    .X(_0942_));
 sky130_fd_sc_hd__xor2_1 _5968_ (.A(_0791_),
    .B(_0794_),
    .X(_0943_));
 sky130_fd_sc_hd__xnor2_1 _5969_ (.A(_0796_),
    .B(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__or2_1 _5970_ (.A(_0942_),
    .B(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__nand2_1 _5971_ (.A(net11),
    .B(net63),
    .Y(_0947_));
 sky130_fd_sc_hd__a21bo_1 _5972_ (.A1(_0942_),
    .A2(_0944_),
    .B1_N(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__a31o_1 _5973_ (.A1(_0811_),
    .A2(_0945_),
    .A3(_0948_),
    .B1(_0812_),
    .X(_0949_));
 sky130_fd_sc_hd__xor2_1 _5974_ (.A(_0652_),
    .B(_0798_),
    .X(_0950_));
 sky130_fd_sc_hd__xnor2_2 _5975_ (.A(_0800_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__nor2_1 _5976_ (.A(_0949_),
    .B(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__and2_1 _5977_ (.A(_0949_),
    .B(_0951_),
    .X(_0953_));
 sky130_fd_sc_hd__and2_1 _5978_ (.A(net14),
    .B(net63),
    .X(_0954_));
 sky130_fd_sc_hd__a21oi_1 _5979_ (.A1(_0949_),
    .A2(_0951_),
    .B1(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__o211a_1 _5980_ (.A1(_0949_),
    .A2(_0951_),
    .B1(net14),
    .C1(net63),
    .X(_0956_));
 sky130_fd_sc_hd__o31a_1 _5981_ (.A1(_0805_),
    .A2(_0953_),
    .A3(_0956_),
    .B1(_0807_),
    .X(_0958_));
 sky130_fd_sc_hd__a31o_1 _5982_ (.A1(_0648_),
    .A2(_0799_),
    .A3(_0801_),
    .B1(_0647_),
    .X(_0959_));
 sky130_fd_sc_hd__nand2b_1 _5983_ (.A_N(_0958_),
    .B(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__and2_1 _5984_ (.A(net63),
    .B(_1716_),
    .X(_0961_));
 sky130_fd_sc_hd__o2bb2a_1 _5985_ (.A1_N(_0960_),
    .A2_N(_0961_),
    .B1(_0044_),
    .B2(_1727_),
    .X(_0962_));
 sky130_fd_sc_hd__and3_1 _5986_ (.A(net64),
    .B(_0960_),
    .C(_0961_),
    .X(_0963_));
 sky130_fd_sc_hd__nor2_1 _5987_ (.A(_0962_),
    .B(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__xnor2_1 _5988_ (.A(_0958_),
    .B(_0959_),
    .Y(_0965_));
 sky130_fd_sc_hd__xnor2_1 _5989_ (.A(_0961_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__nand2_1 _5990_ (.A(net14),
    .B(net64),
    .Y(_0967_));
 sky130_fd_sc_hd__a211o_1 _5991_ (.A1(_0806_),
    .A2(_0807_),
    .B1(_0952_),
    .C1(_0955_),
    .X(_0969_));
 sky130_fd_sc_hd__o211ai_2 _5992_ (.A1(_0952_),
    .A2(_0955_),
    .B1(_0806_),
    .C1(_0807_),
    .Y(_0970_));
 sky130_fd_sc_hd__and3_1 _5993_ (.A(_0967_),
    .B(_0969_),
    .C(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__nand3_1 _5994_ (.A(_0967_),
    .B(_0969_),
    .C(_0970_),
    .Y(_0972_));
 sky130_fd_sc_hd__a21o_1 _5995_ (.A1(_0969_),
    .A2(_0970_),
    .B1(_0967_),
    .X(_0973_));
 sky130_fd_sc_hd__and2_1 _5996_ (.A(net11),
    .B(net64),
    .X(_0974_));
 sky130_fd_sc_hd__a22o_1 _5997_ (.A1(_0811_),
    .A2(_0813_),
    .B1(_0945_),
    .B2(_0948_),
    .X(_0975_));
 sky130_fd_sc_hd__nand4_1 _5998_ (.A(_0811_),
    .B(_0813_),
    .C(_0945_),
    .D(_0948_),
    .Y(_0976_));
 sky130_fd_sc_hd__a21oi_1 _5999_ (.A1(_0975_),
    .A2(_0976_),
    .B1(_0974_),
    .Y(_0977_));
 sky130_fd_sc_hd__a21o_1 _6000_ (.A1(_0975_),
    .A2(_0976_),
    .B1(_0974_),
    .X(_0978_));
 sky130_fd_sc_hd__and3_1 _6001_ (.A(_0974_),
    .B(_0975_),
    .C(_0976_),
    .X(_0980_));
 sky130_fd_sc_hd__a2bb2o_1 _6002_ (.A1_N(_0818_),
    .A2_N(_0820_),
    .B1(_0939_),
    .B2(_0941_),
    .X(_0981_));
 sky130_fd_sc_hd__or4bb_1 _6003_ (.A(_0818_),
    .B(_0820_),
    .C_N(_0939_),
    .D_N(_0941_),
    .X(_0982_));
 sky130_fd_sc_hd__a22o_1 _6004_ (.A1(net9),
    .A2(net64),
    .B1(_0981_),
    .B2(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__and4_1 _6005_ (.A(net9),
    .B(net64),
    .C(_0981_),
    .D(_0982_),
    .X(_0984_));
 sky130_fd_sc_hd__nand4_1 _6006_ (.A(net9),
    .B(net64),
    .C(_0981_),
    .D(_0982_),
    .Y(_0985_));
 sky130_fd_sc_hd__nand2_1 _6007_ (.A(net7),
    .B(net64),
    .Y(_0986_));
 sky130_fd_sc_hd__xnor2_1 _6008_ (.A(_0821_),
    .B(_0823_),
    .Y(_0987_));
 sky130_fd_sc_hd__o21bai_1 _6009_ (.A1(_0833_),
    .A2(_0934_),
    .B1_N(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__or3b_1 _6010_ (.A(_0833_),
    .B(_0934_),
    .C_N(_0987_),
    .X(_0989_));
 sky130_fd_sc_hd__and3_1 _6011_ (.A(_0986_),
    .B(_0988_),
    .C(_0989_),
    .X(_0991_));
 sky130_fd_sc_hd__a21oi_1 _6012_ (.A1(_0988_),
    .A2(_0989_),
    .B1(_0986_),
    .Y(_0992_));
 sky130_fd_sc_hd__nand2_1 _6013_ (.A(net6),
    .B(net64),
    .Y(_0993_));
 sky130_fd_sc_hd__xnor2_1 _6014_ (.A(_0827_),
    .B(_0831_),
    .Y(_0994_));
 sky130_fd_sc_hd__xnor2_1 _6015_ (.A(_0933_),
    .B(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__or2_1 _6016_ (.A(_0993_),
    .B(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__nand2_1 _6017_ (.A(net5),
    .B(net64),
    .Y(_0997_));
 sky130_fd_sc_hd__xor2_1 _6018_ (.A(_0834_),
    .B(_0837_),
    .X(_0998_));
 sky130_fd_sc_hd__xnor2_1 _6019_ (.A(_0932_),
    .B(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__nand2b_1 _6020_ (.A_N(_0997_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__a21oi_1 _6021_ (.A1(net5),
    .A2(net64),
    .B1(_0999_),
    .Y(_1002_));
 sky130_fd_sc_hd__a22o_1 _6022_ (.A1(_0844_),
    .A2(_0846_),
    .B1(_0852_),
    .B2(_0930_),
    .X(_1003_));
 sky130_fd_sc_hd__nand4_2 _6023_ (.A(_0844_),
    .B(_0846_),
    .C(_0852_),
    .D(_0930_),
    .Y(_1004_));
 sky130_fd_sc_hd__and4_1 _6024_ (.A(net4),
    .B(net64),
    .C(_1003_),
    .D(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__a22oi_2 _6025_ (.A1(net4),
    .A2(net64),
    .B1(_1003_),
    .B2(_1004_),
    .Y(_1006_));
 sky130_fd_sc_hd__a22o_1 _6026_ (.A1(net4),
    .A2(net64),
    .B1(_1003_),
    .B2(_1004_),
    .X(_1007_));
 sky130_fd_sc_hd__nand2_1 _6027_ (.A(net3),
    .B(net64),
    .Y(_1008_));
 sky130_fd_sc_hd__inv_2 _6028_ (.A(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__xnor2_1 _6029_ (.A(_0848_),
    .B(_0851_),
    .Y(_1010_));
 sky130_fd_sc_hd__xnor2_1 _6030_ (.A(_0929_),
    .B(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__and2_1 _6031_ (.A(_1009_),
    .B(_1011_),
    .X(_1013_));
 sky130_fd_sc_hd__nand2_1 _6032_ (.A(net2),
    .B(net64),
    .Y(_1014_));
 sky130_fd_sc_hd__inv_2 _6033_ (.A(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__xor2_1 _6034_ (.A(_0853_),
    .B(_0855_),
    .X(_1016_));
 sky130_fd_sc_hd__xnor2_2 _6035_ (.A(_0928_),
    .B(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__and2_1 _6036_ (.A(_1015_),
    .B(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__nand2_1 _6037_ (.A(net32),
    .B(net64),
    .Y(_1019_));
 sky130_fd_sc_hd__inv_2 _6038_ (.A(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__xor2_1 _6039_ (.A(_0859_),
    .B(_0861_),
    .X(_1021_));
 sky130_fd_sc_hd__xnor2_2 _6040_ (.A(_0927_),
    .B(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__and2_1 _6041_ (.A(_1020_),
    .B(_1022_),
    .X(_1024_));
 sky130_fd_sc_hd__a22o_1 _6042_ (.A1(_0867_),
    .A2(_0870_),
    .B1(_0875_),
    .B2(_0926_),
    .X(_1025_));
 sky130_fd_sc_hd__nand4_1 _6043_ (.A(_0867_),
    .B(_0870_),
    .C(_0875_),
    .D(_0926_),
    .Y(_1026_));
 sky130_fd_sc_hd__and4_1 _6044_ (.A(net31),
    .B(net64),
    .C(_1025_),
    .D(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__a22oi_1 _6045_ (.A1(net31),
    .A2(net64),
    .B1(_1025_),
    .B2(_1026_),
    .Y(_1028_));
 sky130_fd_sc_hd__a22o_1 _6046_ (.A1(net31),
    .A2(net64),
    .B1(_1025_),
    .B2(_1026_),
    .X(_1029_));
 sky130_fd_sc_hd__a2bb2o_1 _6047_ (.A1_N(_0873_),
    .A2_N(_0874_),
    .B1(_0881_),
    .B2(_0925_),
    .X(_1030_));
 sky130_fd_sc_hd__or4bb_2 _6048_ (.A(_0873_),
    .B(_0874_),
    .C_N(_0881_),
    .D_N(_0925_),
    .X(_1031_));
 sky130_fd_sc_hd__and4_1 _6049_ (.A(net30),
    .B(net64),
    .C(_1030_),
    .D(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__a22oi_2 _6050_ (.A1(net30),
    .A2(net64),
    .B1(_1030_),
    .B2(_1031_),
    .Y(_1033_));
 sky130_fd_sc_hd__a22o_1 _6051_ (.A1(net30),
    .A2(net64),
    .B1(_1030_),
    .B2(_1031_),
    .X(_1035_));
 sky130_fd_sc_hd__and2_1 _6052_ (.A(net29),
    .B(net64),
    .X(_1036_));
 sky130_fd_sc_hd__xnor2_1 _6053_ (.A(_0876_),
    .B(_0879_),
    .Y(_1037_));
 sky130_fd_sc_hd__xnor2_2 _6054_ (.A(_0923_),
    .B(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__and2_1 _6055_ (.A(_1036_),
    .B(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__xor2_1 _6056_ (.A(_0882_),
    .B(_0884_),
    .X(_1040_));
 sky130_fd_sc_hd__xnor2_2 _6057_ (.A(_0922_),
    .B(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__and2_1 _6058_ (.A(net28),
    .B(net64),
    .X(_1042_));
 sky130_fd_sc_hd__or2_1 _6059_ (.A(_1041_),
    .B(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__a21o_1 _6060_ (.A1(_0890_),
    .A2(_0892_),
    .B1(_0921_),
    .X(_1044_));
 sky130_fd_sc_hd__nand3_1 _6061_ (.A(_0890_),
    .B(_0892_),
    .C(_0921_),
    .Y(_1046_));
 sky130_fd_sc_hd__a22o_1 _6062_ (.A1(net27),
    .A2(net64),
    .B1(_1044_),
    .B2(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__and4_1 _6063_ (.A(net27),
    .B(net64),
    .C(_1044_),
    .D(_1046_),
    .X(_1048_));
 sky130_fd_sc_hd__nand4_1 _6064_ (.A(net27),
    .B(net64),
    .C(_1044_),
    .D(_1046_),
    .Y(_1049_));
 sky130_fd_sc_hd__nand2_1 _6065_ (.A(net26),
    .B(net64),
    .Y(_1050_));
 sky130_fd_sc_hd__o22ai_2 _6066_ (.A1(_0896_),
    .A2(_0897_),
    .B1(_0904_),
    .B2(_0920_),
    .Y(_1051_));
 sky130_fd_sc_hd__or4_1 _6067_ (.A(_0896_),
    .B(_0897_),
    .C(_0904_),
    .D(_0920_),
    .X(_1052_));
 sky130_fd_sc_hd__and3_1 _6068_ (.A(_1050_),
    .B(_1051_),
    .C(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__nand3_1 _6069_ (.A(_1050_),
    .B(_1051_),
    .C(_1052_),
    .Y(_1054_));
 sky130_fd_sc_hd__a21oi_1 _6070_ (.A1(_1051_),
    .A2(_1052_),
    .B1(_1050_),
    .Y(_1055_));
 sky130_fd_sc_hd__nand2_1 _6071_ (.A(net23),
    .B(net64),
    .Y(_1057_));
 sky130_fd_sc_hd__xnor2_1 _6072_ (.A(_0899_),
    .B(_0903_),
    .Y(_1058_));
 sky130_fd_sc_hd__xnor2_2 _6073_ (.A(_0919_),
    .B(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__a21o_1 _6074_ (.A1(net23),
    .A2(net64),
    .B1(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__nand2_1 _6075_ (.A(net12),
    .B(net64),
    .Y(_1061_));
 sky130_fd_sc_hd__inv_2 _6076_ (.A(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__xor2_1 _6077_ (.A(_0905_),
    .B(_0907_),
    .X(_1063_));
 sky130_fd_sc_hd__xnor2_1 _6078_ (.A(_0918_),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__and2_1 _6079_ (.A(_1062_),
    .B(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__a21oi_1 _6080_ (.A1(_0912_),
    .A2(_0914_),
    .B1(_0917_),
    .Y(_1066_));
 sky130_fd_sc_hd__and3_1 _6081_ (.A(_0912_),
    .B(_0914_),
    .C(_0917_),
    .X(_1068_));
 sky130_fd_sc_hd__o211ai_2 _6082_ (.A1(_1066_),
    .A2(_1068_),
    .B1(net1),
    .C1(net64),
    .Y(_1069_));
 sky130_fd_sc_hd__o21ba_1 _6083_ (.A1(_1062_),
    .A2(_1064_),
    .B1_N(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__nor2_1 _6084_ (.A(_1065_),
    .B(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__a311o_1 _6085_ (.A1(net23),
    .A2(net64),
    .A3(_1059_),
    .B1(_1065_),
    .C1(_1070_),
    .X(_1072_));
 sky130_fd_sc_hd__a31o_1 _6086_ (.A1(_1054_),
    .A2(_1060_),
    .A3(_1072_),
    .B1(_1055_),
    .X(_1073_));
 sky130_fd_sc_hd__a21oi_1 _6087_ (.A1(_1047_),
    .A2(_1073_),
    .B1(_1048_),
    .Y(_1074_));
 sky130_fd_sc_hd__a221o_1 _6088_ (.A1(_1041_),
    .A2(_1042_),
    .B1(_1047_),
    .B2(_1073_),
    .C1(_1048_),
    .X(_1075_));
 sky130_fd_sc_hd__nand2_1 _6089_ (.A(_1043_),
    .B(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__o211a_1 _6090_ (.A1(_1036_),
    .A2(_1038_),
    .B1(_1043_),
    .C1(_1075_),
    .X(_1077_));
 sky130_fd_sc_hd__o31ai_1 _6091_ (.A1(_1032_),
    .A2(_1039_),
    .A3(_1077_),
    .B1(_1035_),
    .Y(_1079_));
 sky130_fd_sc_hd__o31a_1 _6092_ (.A1(_1032_),
    .A2(_1039_),
    .A3(_1077_),
    .B1(_1035_),
    .X(_1080_));
 sky130_fd_sc_hd__o21a_1 _6093_ (.A1(_1027_),
    .A2(_1080_),
    .B1(_1029_),
    .X(_1081_));
 sky130_fd_sc_hd__o221a_1 _6094_ (.A1(_1020_),
    .A2(_1022_),
    .B1(_1027_),
    .B2(_1080_),
    .C1(_1029_),
    .X(_1082_));
 sky130_fd_sc_hd__or2_1 _6095_ (.A(_1024_),
    .B(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__o22a_1 _6096_ (.A1(_1015_),
    .A2(_1017_),
    .B1(_1024_),
    .B2(_1082_),
    .X(_1084_));
 sky130_fd_sc_hd__nor2_1 _6097_ (.A(_1018_),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__o22a_1 _6098_ (.A1(_1009_),
    .A2(_1011_),
    .B1(_1018_),
    .B2(_1084_),
    .X(_1086_));
 sky130_fd_sc_hd__o31ai_2 _6099_ (.A1(_1005_),
    .A2(_1013_),
    .A3(_1086_),
    .B1(_1007_),
    .Y(_1087_));
 sky130_fd_sc_hd__a21oi_1 _6100_ (.A1(_1000_),
    .A2(_1087_),
    .B1(_1002_),
    .Y(_1088_));
 sky130_fd_sc_hd__a221o_1 _6101_ (.A1(_0993_),
    .A2(_0995_),
    .B1(_1000_),
    .B2(_1087_),
    .C1(_1002_),
    .X(_1090_));
 sky130_fd_sc_hd__nand2_1 _6102_ (.A(_0996_),
    .B(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__and3b_1 _6103_ (.A_N(_0992_),
    .B(_0996_),
    .C(_1090_),
    .X(_1092_));
 sky130_fd_sc_hd__a21oi_1 _6104_ (.A1(_0996_),
    .A2(_1090_),
    .B1(_0991_),
    .Y(_1093_));
 sky130_fd_sc_hd__xor2_1 _6105_ (.A(_0936_),
    .B(_0938_),
    .X(_1094_));
 sky130_fd_sc_hd__xor2_1 _6106_ (.A(_0940_),
    .B(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__xnor2_1 _6107_ (.A(_0940_),
    .B(_1094_),
    .Y(_1096_));
 sky130_fd_sc_hd__o21a_1 _6108_ (.A1(_0991_),
    .A2(_1092_),
    .B1(_1095_),
    .X(_1097_));
 sky130_fd_sc_hd__o21a_1 _6109_ (.A1(_0992_),
    .A2(_1093_),
    .B1(_1096_),
    .X(_1098_));
 sky130_fd_sc_hd__nand2_1 _6110_ (.A(net8),
    .B(net64),
    .Y(_1099_));
 sky130_fd_sc_hd__o31a_1 _6111_ (.A1(_0991_),
    .A2(_1092_),
    .A3(_1095_),
    .B1(_1099_),
    .X(_1101_));
 sky130_fd_sc_hd__o311a_1 _6112_ (.A1(_0992_),
    .A2(_1093_),
    .A3(_1096_),
    .B1(net64),
    .C1(net8),
    .X(_1102_));
 sky130_fd_sc_hd__o31a_1 _6113_ (.A1(_0984_),
    .A2(_1098_),
    .A3(_1102_),
    .B1(_0983_),
    .X(_1103_));
 sky130_fd_sc_hd__xor2_1 _6114_ (.A(_0942_),
    .B(_0944_),
    .X(_1104_));
 sky130_fd_sc_hd__xnor2_1 _6115_ (.A(_0947_),
    .B(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__or2_1 _6116_ (.A(_1103_),
    .B(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__and2_1 _6117_ (.A(net10),
    .B(net64),
    .X(_1107_));
 sky130_fd_sc_hd__a21o_1 _6118_ (.A1(_1103_),
    .A2(_1105_),
    .B1(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__a31o_1 _6119_ (.A1(_0978_),
    .A2(_1106_),
    .A3(_1108_),
    .B1(_0980_),
    .X(_1109_));
 sky130_fd_sc_hd__xnor2_1 _6120_ (.A(_0949_),
    .B(_0951_),
    .Y(_1110_));
 sky130_fd_sc_hd__xnor2_2 _6121_ (.A(_0954_),
    .B(_1110_),
    .Y(_1112_));
 sky130_fd_sc_hd__or2_1 _6122_ (.A(_1109_),
    .B(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__nand2_1 _6123_ (.A(_1109_),
    .B(_1112_),
    .Y(_1114_));
 sky130_fd_sc_hd__nand2_1 _6124_ (.A(net13),
    .B(net64),
    .Y(_1115_));
 sky130_fd_sc_hd__a21bo_1 _6125_ (.A1(_1109_),
    .A2(_1112_),
    .B1_N(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__o211ai_1 _6126_ (.A1(_1109_),
    .A2(_1112_),
    .B1(net13),
    .C1(net64),
    .Y(_1117_));
 sky130_fd_sc_hd__a31o_1 _6127_ (.A1(_0973_),
    .A2(_1114_),
    .A3(_1117_),
    .B1(_0971_),
    .X(_1118_));
 sky130_fd_sc_hd__or2_1 _6128_ (.A(_0966_),
    .B(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__nand2_1 _6129_ (.A(net15),
    .B(net64),
    .Y(_1120_));
 sky130_fd_sc_hd__a21o_1 _6130_ (.A1(_0966_),
    .A2(_1118_),
    .B1(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__a21o_1 _6131_ (.A1(_1119_),
    .A2(_1121_),
    .B1(_0964_),
    .X(_1123_));
 sky130_fd_sc_hd__nand3_1 _6132_ (.A(_0964_),
    .B(_1119_),
    .C(_1121_),
    .Y(_1124_));
 sky130_fd_sc_hd__and3_1 _6133_ (.A(_3985_),
    .B(_1123_),
    .C(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__nand3_2 _6134_ (.A(_3985_),
    .B(_1123_),
    .C(_1124_),
    .Y(_1126_));
 sky130_fd_sc_hd__a21oi_2 _6135_ (.A1(_1123_),
    .A2(_1124_),
    .B1(_3985_),
    .Y(_1127_));
 sky130_fd_sc_hd__and2_1 _6136_ (.A(net13),
    .B(net34),
    .X(_1128_));
 sky130_fd_sc_hd__a22o_1 _6137_ (.A1(_0972_),
    .A2(_0973_),
    .B1(_1113_),
    .B2(_1116_),
    .X(_1129_));
 sky130_fd_sc_hd__nand4_1 _6138_ (.A(_0972_),
    .B(_0973_),
    .C(_1113_),
    .D(_1116_),
    .Y(_1130_));
 sky130_fd_sc_hd__and3_1 _6139_ (.A(_1128_),
    .B(_1129_),
    .C(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__a21oi_1 _6140_ (.A1(_1129_),
    .A2(_1130_),
    .B1(_1128_),
    .Y(_1132_));
 sky130_fd_sc_hd__a21o_1 _6141_ (.A1(_1129_),
    .A2(_1130_),
    .B1(_1128_),
    .X(_1134_));
 sky130_fd_sc_hd__xor2_1 _6142_ (.A(_1109_),
    .B(_1112_),
    .X(_1135_));
 sky130_fd_sc_hd__xnor2_1 _6143_ (.A(_1115_),
    .B(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__and2_1 _6144_ (.A(net10),
    .B(net34),
    .X(_1137_));
 sky130_fd_sc_hd__a2bb2o_1 _6145_ (.A1_N(_0977_),
    .A2_N(_0980_),
    .B1(_1106_),
    .B2(_1108_),
    .X(_1138_));
 sky130_fd_sc_hd__or4bb_1 _6146_ (.A(_0977_),
    .B(_0980_),
    .C_N(_1106_),
    .D_N(_1108_),
    .X(_1139_));
 sky130_fd_sc_hd__a21o_1 _6147_ (.A1(_1138_),
    .A2(_1139_),
    .B1(_1137_),
    .X(_1140_));
 sky130_fd_sc_hd__and3_1 _6148_ (.A(_1137_),
    .B(_1138_),
    .C(_1139_),
    .X(_1141_));
 sky130_fd_sc_hd__nand3_1 _6149_ (.A(_1137_),
    .B(_1138_),
    .C(_1139_),
    .Y(_1142_));
 sky130_fd_sc_hd__and2_1 _6150_ (.A(net8),
    .B(net34),
    .X(_1143_));
 sky130_fd_sc_hd__o2bb2a_1 _6151_ (.A1_N(_0983_),
    .A2_N(_0985_),
    .B1(_1098_),
    .B2(_1102_),
    .X(_1145_));
 sky130_fd_sc_hd__o211a_1 _6152_ (.A1(_1097_),
    .A2(_1101_),
    .B1(_0983_),
    .C1(_0985_),
    .X(_1146_));
 sky130_fd_sc_hd__or3_1 _6153_ (.A(_1143_),
    .B(_1145_),
    .C(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__o21a_1 _6154_ (.A1(_1145_),
    .A2(_1146_),
    .B1(_1143_),
    .X(_1148_));
 sky130_fd_sc_hd__o21ai_1 _6155_ (.A1(_1145_),
    .A2(_1146_),
    .B1(_1143_),
    .Y(_1149_));
 sky130_fd_sc_hd__or3_1 _6156_ (.A(_1097_),
    .B(_1098_),
    .C(_1099_),
    .X(_1150_));
 sky130_fd_sc_hd__o21ai_1 _6157_ (.A1(_1097_),
    .A2(_1098_),
    .B1(_1099_),
    .Y(_1151_));
 sky130_fd_sc_hd__nand2_1 _6158_ (.A(net6),
    .B(net34),
    .Y(_1152_));
 sky130_fd_sc_hd__or2_1 _6159_ (.A(_0991_),
    .B(_0992_),
    .X(_1153_));
 sky130_fd_sc_hd__xnor2_1 _6160_ (.A(_1091_),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__nand2b_1 _6161_ (.A_N(_1154_),
    .B(_1152_),
    .Y(_1156_));
 sky130_fd_sc_hd__and2_1 _6162_ (.A(net5),
    .B(net34),
    .X(_1157_));
 sky130_fd_sc_hd__xnor2_1 _6163_ (.A(_0993_),
    .B(_0995_),
    .Y(_1158_));
 sky130_fd_sc_hd__xnor2_1 _6164_ (.A(_1088_),
    .B(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__or2_1 _6165_ (.A(_1157_),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__nand2_1 _6166_ (.A(net4),
    .B(net34),
    .Y(_1161_));
 sky130_fd_sc_hd__xnor2_1 _6167_ (.A(_0997_),
    .B(_0999_),
    .Y(_1162_));
 sky130_fd_sc_hd__xnor2_1 _6168_ (.A(_1087_),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__and3_1 _6169_ (.A(net4),
    .B(net34),
    .C(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__a21o_1 _6170_ (.A1(net4),
    .A2(net34),
    .B1(_1163_),
    .X(_1165_));
 sky130_fd_sc_hd__nand2_1 _6171_ (.A(net3),
    .B(net34),
    .Y(_1167_));
 sky130_fd_sc_hd__o22ai_2 _6172_ (.A1(_1005_),
    .A2(_1006_),
    .B1(_1013_),
    .B2(_1086_),
    .Y(_1168_));
 sky130_fd_sc_hd__or4_1 _6173_ (.A(_1005_),
    .B(_1006_),
    .C(_1013_),
    .D(_1086_),
    .X(_1169_));
 sky130_fd_sc_hd__a21oi_1 _6174_ (.A1(_1168_),
    .A2(_1169_),
    .B1(_1167_),
    .Y(_1170_));
 sky130_fd_sc_hd__a21o_1 _6175_ (.A1(_1168_),
    .A2(_1169_),
    .B1(_1167_),
    .X(_1171_));
 sky130_fd_sc_hd__and3_1 _6176_ (.A(_1167_),
    .B(_1168_),
    .C(_1169_),
    .X(_1172_));
 sky130_fd_sc_hd__nand2_1 _6177_ (.A(net2),
    .B(net34),
    .Y(_1173_));
 sky130_fd_sc_hd__inv_2 _6178_ (.A(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__xnor2_1 _6179_ (.A(_1008_),
    .B(_1011_),
    .Y(_1175_));
 sky130_fd_sc_hd__xnor2_2 _6180_ (.A(_1085_),
    .B(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__nand2_1 _6181_ (.A(_1174_),
    .B(_1176_),
    .Y(_1178_));
 sky130_fd_sc_hd__nand2_1 _6182_ (.A(net32),
    .B(net34),
    .Y(_1179_));
 sky130_fd_sc_hd__xnor2_1 _6183_ (.A(_1015_),
    .B(_1017_),
    .Y(_1180_));
 sky130_fd_sc_hd__xnor2_1 _6184_ (.A(_1083_),
    .B(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__and3_1 _6185_ (.A(net32),
    .B(net34),
    .C(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__nand2b_1 _6186_ (.A_N(_1181_),
    .B(_1179_),
    .Y(_1183_));
 sky130_fd_sc_hd__nand2_1 _6187_ (.A(net31),
    .B(net34),
    .Y(_1184_));
 sky130_fd_sc_hd__xnor2_1 _6188_ (.A(_1020_),
    .B(_1022_),
    .Y(_1185_));
 sky130_fd_sc_hd__xnor2_1 _6189_ (.A(_1081_),
    .B(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__and3_1 _6190_ (.A(net31),
    .B(net34),
    .C(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__nand2b_1 _6191_ (.A_N(_1186_),
    .B(_1184_),
    .Y(_1189_));
 sky130_fd_sc_hd__o21ai_1 _6192_ (.A1(_1027_),
    .A2(_1028_),
    .B1(_1079_),
    .Y(_1190_));
 sky130_fd_sc_hd__or3_1 _6193_ (.A(_1027_),
    .B(_1028_),
    .C(_1079_),
    .X(_1191_));
 sky130_fd_sc_hd__nand4_1 _6194_ (.A(net30),
    .B(net34),
    .C(_1190_),
    .D(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__a22o_1 _6195_ (.A1(net30),
    .A2(net34),
    .B1(_1190_),
    .B2(_1191_),
    .X(_1193_));
 sky130_fd_sc_hd__nand2_1 _6196_ (.A(net29),
    .B(net34),
    .Y(_1194_));
 sky130_fd_sc_hd__o22ai_2 _6197_ (.A1(_1032_),
    .A2(_1033_),
    .B1(_1039_),
    .B2(_1077_),
    .Y(_1195_));
 sky130_fd_sc_hd__or4_1 _6198_ (.A(_1032_),
    .B(_1033_),
    .C(_1039_),
    .D(_1077_),
    .X(_1196_));
 sky130_fd_sc_hd__nand3_2 _6199_ (.A(_1194_),
    .B(_1195_),
    .C(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__a21oi_1 _6200_ (.A1(_1195_),
    .A2(_1196_),
    .B1(_1194_),
    .Y(_1198_));
 sky130_fd_sc_hd__a21o_1 _6201_ (.A1(_1195_),
    .A2(_1196_),
    .B1(_1194_),
    .X(_1200_));
 sky130_fd_sc_hd__nand2_2 _6202_ (.A(net28),
    .B(net34),
    .Y(_1201_));
 sky130_fd_sc_hd__xor2_1 _6203_ (.A(_1036_),
    .B(_1038_),
    .X(_1202_));
 sky130_fd_sc_hd__xor2_2 _6204_ (.A(_1076_),
    .B(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__nor2_1 _6205_ (.A(_1201_),
    .B(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__nand2_1 _6206_ (.A(net27),
    .B(net34),
    .Y(_1205_));
 sky130_fd_sc_hd__xor2_1 _6207_ (.A(_1041_),
    .B(_1042_),
    .X(_1206_));
 sky130_fd_sc_hd__xnor2_2 _6208_ (.A(_1074_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__nand2b_1 _6209_ (.A_N(_1205_),
    .B(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__a21oi_2 _6210_ (.A1(net27),
    .A2(net34),
    .B1(_1207_),
    .Y(_1209_));
 sky130_fd_sc_hd__a21o_1 _6211_ (.A1(_1047_),
    .A2(_1049_),
    .B1(_1073_),
    .X(_1211_));
 sky130_fd_sc_hd__nand3_1 _6212_ (.A(_1047_),
    .B(_1049_),
    .C(_1073_),
    .Y(_1212_));
 sky130_fd_sc_hd__and4_1 _6213_ (.A(net26),
    .B(net34),
    .C(_1211_),
    .D(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__nand4_1 _6214_ (.A(net26),
    .B(net34),
    .C(_1211_),
    .D(_1212_),
    .Y(_1214_));
 sky130_fd_sc_hd__a22oi_2 _6215_ (.A1(net26),
    .A2(net34),
    .B1(_1211_),
    .B2(_1212_),
    .Y(_1215_));
 sky130_fd_sc_hd__nand2_1 _6216_ (.A(net23),
    .B(net34),
    .Y(_1216_));
 sky130_fd_sc_hd__o211ai_1 _6217_ (.A1(_1053_),
    .A2(_1055_),
    .B1(_1060_),
    .C1(_1072_),
    .Y(_1217_));
 sky130_fd_sc_hd__a211o_1 _6218_ (.A1(_1060_),
    .A2(_1072_),
    .B1(_1053_),
    .C1(_1055_),
    .X(_1218_));
 sky130_fd_sc_hd__and3_1 _6219_ (.A(_1216_),
    .B(_1217_),
    .C(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__a21oi_2 _6220_ (.A1(_1217_),
    .A2(_1218_),
    .B1(_1216_),
    .Y(_1220_));
 sky130_fd_sc_hd__xnor2_1 _6221_ (.A(_1057_),
    .B(_1059_),
    .Y(_1222_));
 sky130_fd_sc_hd__xnor2_1 _6222_ (.A(_1071_),
    .B(_1222_),
    .Y(_1223_));
 sky130_fd_sc_hd__and2_1 _6223_ (.A(net12),
    .B(net34),
    .X(_1224_));
 sky130_fd_sc_hd__nand2_1 _6224_ (.A(_1223_),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__or2_1 _6225_ (.A(_1223_),
    .B(_1224_),
    .X(_1226_));
 sky130_fd_sc_hd__xnor2_1 _6226_ (.A(_1062_),
    .B(_1064_),
    .Y(_1227_));
 sky130_fd_sc_hd__o211a_1 _6227_ (.A1(_1069_),
    .A2(_1227_),
    .B1(net1),
    .C1(net34),
    .X(_1228_));
 sky130_fd_sc_hd__a21bo_1 _6228_ (.A1(_1069_),
    .A2(_1227_),
    .B1_N(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__o21bai_2 _6229_ (.A1(_1223_),
    .A2(_1224_),
    .B1_N(_1229_),
    .Y(_1230_));
 sky130_fd_sc_hd__and3b_1 _6230_ (.A_N(_1220_),
    .B(_1225_),
    .C(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__a21oi_1 _6231_ (.A1(_1225_),
    .A2(_1230_),
    .B1(_1219_),
    .Y(_1233_));
 sky130_fd_sc_hd__o31a_2 _6232_ (.A1(_1215_),
    .A2(_1219_),
    .A3(_1231_),
    .B1(_1214_),
    .X(_1234_));
 sky130_fd_sc_hd__a21o_1 _6233_ (.A1(_1208_),
    .A2(_1234_),
    .B1(_1209_),
    .X(_1235_));
 sky130_fd_sc_hd__a221oi_4 _6234_ (.A1(_1201_),
    .A2(_1203_),
    .B1(_1208_),
    .B2(_1234_),
    .C1(_1209_),
    .Y(_1236_));
 sky130_fd_sc_hd__o31ai_2 _6235_ (.A1(_1198_),
    .A2(_1204_),
    .A3(_1236_),
    .B1(_1197_),
    .Y(_1237_));
 sky130_fd_sc_hd__a21boi_1 _6236_ (.A1(_1192_),
    .A2(_1237_),
    .B1_N(_1193_),
    .Y(_1238_));
 sky130_fd_sc_hd__o21a_1 _6237_ (.A1(_1187_),
    .A2(_1238_),
    .B1(_1189_),
    .X(_1239_));
 sky130_fd_sc_hd__o21ai_1 _6238_ (.A1(_1182_),
    .A2(_1239_),
    .B1(_1183_),
    .Y(_1240_));
 sky130_fd_sc_hd__o221ai_4 _6239_ (.A1(_1174_),
    .A2(_1176_),
    .B1(_1182_),
    .B2(_1239_),
    .C1(_1183_),
    .Y(_1241_));
 sky130_fd_sc_hd__a31oi_2 _6240_ (.A1(_1171_),
    .A2(_1178_),
    .A3(_1241_),
    .B1(_1172_),
    .Y(_1242_));
 sky130_fd_sc_hd__a21o_1 _6241_ (.A1(_1165_),
    .A2(_1242_),
    .B1(_1164_),
    .X(_1244_));
 sky130_fd_sc_hd__a221o_1 _6242_ (.A1(_1157_),
    .A2(_1159_),
    .B1(_1165_),
    .B2(_1242_),
    .C1(_1164_),
    .X(_1245_));
 sky130_fd_sc_hd__nand2_1 _6243_ (.A(_1160_),
    .B(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__a32o_1 _6244_ (.A1(net6),
    .A2(net34),
    .A3(_1154_),
    .B1(_1160_),
    .B2(_1245_),
    .X(_1247_));
 sky130_fd_sc_hd__a22o_1 _6245_ (.A1(_1150_),
    .A2(_1151_),
    .B1(_1156_),
    .B2(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__nand4_1 _6246_ (.A(_1150_),
    .B(_1151_),
    .C(_1156_),
    .D(_1247_),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_1 _6247_ (.A(net7),
    .B(net34),
    .Y(_1250_));
 sky130_fd_sc_hd__inv_2 _6248_ (.A(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__a41o_1 _6249_ (.A1(_1150_),
    .A2(_1151_),
    .A3(_1156_),
    .A4(_1247_),
    .B1(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__a31o_1 _6250_ (.A1(_1147_),
    .A2(_1248_),
    .A3(_1252_),
    .B1(_1148_),
    .X(_1253_));
 sky130_fd_sc_hd__xor2_1 _6251_ (.A(_1103_),
    .B(_1105_),
    .X(_1255_));
 sky130_fd_sc_hd__xor2_1 _6252_ (.A(_1107_),
    .B(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__or2_1 _6253_ (.A(_1253_),
    .B(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__nand2_1 _6254_ (.A(net9),
    .B(net34),
    .Y(_1258_));
 sky130_fd_sc_hd__a21bo_1 _6255_ (.A1(_1253_),
    .A2(_1256_),
    .B1_N(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__a31o_1 _6256_ (.A1(_1140_),
    .A2(_1257_),
    .A3(_1259_),
    .B1(_1141_),
    .X(_1260_));
 sky130_fd_sc_hd__or2_1 _6257_ (.A(_1136_),
    .B(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__nand2_1 _6258_ (.A(net11),
    .B(net34),
    .Y(_1262_));
 sky130_fd_sc_hd__a21bo_1 _6259_ (.A1(_1136_),
    .A2(_1260_),
    .B1_N(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__a31o_1 _6260_ (.A1(_1134_),
    .A2(_1261_),
    .A3(_1263_),
    .B1(_1131_),
    .X(_1264_));
 sky130_fd_sc_hd__xor2_1 _6261_ (.A(_0966_),
    .B(_1118_),
    .X(_1266_));
 sky130_fd_sc_hd__xnor2_1 _6262_ (.A(_1120_),
    .B(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__or2_1 _6263_ (.A(_1264_),
    .B(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__nand2_1 _6264_ (.A(net14),
    .B(net34),
    .Y(_1269_));
 sky130_fd_sc_hd__a21bo_1 _6265_ (.A1(_1264_),
    .A2(_1267_),
    .B1_N(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__and2_1 _6266_ (.A(_1268_),
    .B(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__a21oi_1 _6267_ (.A1(_1268_),
    .A2(_1270_),
    .B1(_1127_),
    .Y(_1272_));
 sky130_fd_sc_hd__a31oi_2 _6268_ (.A1(_1126_),
    .A2(_1268_),
    .A3(_1270_),
    .B1(_1127_),
    .Y(_1273_));
 sky130_fd_sc_hd__a21oi_1 _6269_ (.A1(_1119_),
    .A2(_1121_),
    .B1(_0962_),
    .Y(_1274_));
 sky130_fd_sc_hd__or2_1 _6270_ (.A(_0963_),
    .B(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__a211o_1 _6271_ (.A1(_1126_),
    .A2(_1271_),
    .B1(_1275_),
    .C1(_1127_),
    .X(_1277_));
 sky130_fd_sc_hd__a31o_1 _6272_ (.A1(net34),
    .A2(_1716_),
    .A3(_1277_),
    .B1(_3983_),
    .X(_1278_));
 sky130_fd_sc_hd__or3b_1 _6273_ (.A(_0055_),
    .B(_3984_),
    .C_N(_1277_),
    .X(_1279_));
 sky130_fd_sc_hd__and2_1 _6274_ (.A(_1278_),
    .B(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__xor2_1 _6275_ (.A(_1273_),
    .B(_1275_),
    .X(_1281_));
 sky130_fd_sc_hd__xnor2_1 _6276_ (.A(_3984_),
    .B(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__and2_1 _6277_ (.A(net14),
    .B(net35),
    .X(_1283_));
 sky130_fd_sc_hd__or2_1 _6278_ (.A(_1125_),
    .B(_1127_),
    .X(_1284_));
 sky130_fd_sc_hd__and3_1 _6279_ (.A(_1127_),
    .B(_1268_),
    .C(_1270_),
    .X(_1285_));
 sky130_fd_sc_hd__a221oi_1 _6280_ (.A1(_1126_),
    .A2(_1272_),
    .B1(_1284_),
    .B2(_1271_),
    .C1(_1283_),
    .Y(_1286_));
 sky130_fd_sc_hd__a221o_1 _6281_ (.A1(_1126_),
    .A2(_1272_),
    .B1(_1284_),
    .B2(_1271_),
    .C1(_1283_),
    .X(_1288_));
 sky130_fd_sc_hd__o221a_1 _6282_ (.A1(_1126_),
    .A2(_1271_),
    .B1(_1273_),
    .B2(_1285_),
    .C1(_1283_),
    .X(_1289_));
 sky130_fd_sc_hd__nand2_1 _6283_ (.A(net11),
    .B(net35),
    .Y(_1290_));
 sky130_fd_sc_hd__o211ai_2 _6284_ (.A1(_1131_),
    .A2(_1132_),
    .B1(_1261_),
    .C1(_1263_),
    .Y(_1291_));
 sky130_fd_sc_hd__a211o_1 _6285_ (.A1(_1261_),
    .A2(_1263_),
    .B1(_1131_),
    .C1(_1132_),
    .X(_1292_));
 sky130_fd_sc_hd__a21oi_1 _6286_ (.A1(_1291_),
    .A2(_1292_),
    .B1(_1290_),
    .Y(_1293_));
 sky130_fd_sc_hd__a21o_1 _6287_ (.A1(_1291_),
    .A2(_1292_),
    .B1(_1290_),
    .X(_1294_));
 sky130_fd_sc_hd__and3_1 _6288_ (.A(_1290_),
    .B(_1291_),
    .C(_1292_),
    .X(_1295_));
 sky130_fd_sc_hd__a22o_1 _6289_ (.A1(_1140_),
    .A2(_1142_),
    .B1(_1257_),
    .B2(_1259_),
    .X(_1296_));
 sky130_fd_sc_hd__nand4_1 _6290_ (.A(_1140_),
    .B(_1142_),
    .C(_1257_),
    .D(_1259_),
    .Y(_1297_));
 sky130_fd_sc_hd__and4_1 _6291_ (.A(net9),
    .B(net35),
    .C(_1296_),
    .D(_1297_),
    .X(_1299_));
 sky130_fd_sc_hd__nand4_1 _6292_ (.A(net9),
    .B(net35),
    .C(_1296_),
    .D(_1297_),
    .Y(_1300_));
 sky130_fd_sc_hd__a22o_1 _6293_ (.A1(net9),
    .A2(net35),
    .B1(_1296_),
    .B2(_1297_),
    .X(_1301_));
 sky130_fd_sc_hd__and2_1 _6294_ (.A(net7),
    .B(net35),
    .X(_1302_));
 sky130_fd_sc_hd__a22o_1 _6295_ (.A1(_1147_),
    .A2(_1149_),
    .B1(_1248_),
    .B2(_1252_),
    .X(_1303_));
 sky130_fd_sc_hd__nand4_2 _6296_ (.A(_1147_),
    .B(_1149_),
    .C(_1248_),
    .D(_1252_),
    .Y(_1304_));
 sky130_fd_sc_hd__a21oi_2 _6297_ (.A1(_1303_),
    .A2(_1304_),
    .B1(_1302_),
    .Y(_1305_));
 sky130_fd_sc_hd__a21o_1 _6298_ (.A1(_1303_),
    .A2(_1304_),
    .B1(_1302_),
    .X(_1306_));
 sky130_fd_sc_hd__and3_1 _6299_ (.A(_1302_),
    .B(_1303_),
    .C(_1304_),
    .X(_1307_));
 sky130_fd_sc_hd__and3_1 _6300_ (.A(_1248_),
    .B(_1249_),
    .C(_1250_),
    .X(_1308_));
 sky130_fd_sc_hd__a21oi_2 _6301_ (.A1(_1248_),
    .A2(_1249_),
    .B1(_1250_),
    .Y(_1310_));
 sky130_fd_sc_hd__and2_1 _6302_ (.A(net5),
    .B(net35),
    .X(_1311_));
 sky130_fd_sc_hd__xnor2_1 _6303_ (.A(_1152_),
    .B(_1154_),
    .Y(_1312_));
 sky130_fd_sc_hd__xnor2_1 _6304_ (.A(_1246_),
    .B(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__and2_1 _6305_ (.A(_1311_),
    .B(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__nand2_1 _6306_ (.A(net4),
    .B(net35),
    .Y(_1315_));
 sky130_fd_sc_hd__xnor2_1 _6307_ (.A(_1157_),
    .B(_1159_),
    .Y(_1316_));
 sky130_fd_sc_hd__xnor2_1 _6308_ (.A(_1244_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__nand2b_1 _6309_ (.A_N(_1317_),
    .B(_1315_),
    .Y(_1318_));
 sky130_fd_sc_hd__and3_1 _6310_ (.A(net4),
    .B(net35),
    .C(_1317_),
    .X(_1319_));
 sky130_fd_sc_hd__nand2_1 _6311_ (.A(net3),
    .B(net35),
    .Y(_1321_));
 sky130_fd_sc_hd__xor2_1 _6312_ (.A(_1161_),
    .B(_1163_),
    .X(_1322_));
 sky130_fd_sc_hd__xnor2_1 _6313_ (.A(_1242_),
    .B(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__a21o_1 _6314_ (.A1(net3),
    .A2(net35),
    .B1(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__and3_1 _6315_ (.A(net3),
    .B(net35),
    .C(_1323_),
    .X(_1325_));
 sky130_fd_sc_hd__and2_1 _6316_ (.A(net2),
    .B(net35),
    .X(_1326_));
 sky130_fd_sc_hd__o211ai_2 _6317_ (.A1(_1170_),
    .A2(_1172_),
    .B1(_1178_),
    .C1(_1241_),
    .Y(_1327_));
 sky130_fd_sc_hd__a211o_1 _6318_ (.A1(_1178_),
    .A2(_1241_),
    .B1(_1170_),
    .C1(_1172_),
    .X(_1328_));
 sky130_fd_sc_hd__a21o_1 _6319_ (.A1(_1327_),
    .A2(_1328_),
    .B1(_1326_),
    .X(_1329_));
 sky130_fd_sc_hd__and3_1 _6320_ (.A(_1326_),
    .B(_1327_),
    .C(_1328_),
    .X(_1330_));
 sky130_fd_sc_hd__nand3_1 _6321_ (.A(_1326_),
    .B(_1327_),
    .C(_1328_),
    .Y(_1332_));
 sky130_fd_sc_hd__and2_1 _6322_ (.A(net32),
    .B(net35),
    .X(_1333_));
 sky130_fd_sc_hd__xnor2_1 _6323_ (.A(_1173_),
    .B(_1176_),
    .Y(_1334_));
 sky130_fd_sc_hd__xnor2_2 _6324_ (.A(_1240_),
    .B(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__and2_1 _6325_ (.A(_1333_),
    .B(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__or2_1 _6326_ (.A(_1333_),
    .B(_1335_),
    .X(_1337_));
 sky130_fd_sc_hd__and2_1 _6327_ (.A(net31),
    .B(net35),
    .X(_1338_));
 sky130_fd_sc_hd__xor2_1 _6328_ (.A(_1179_),
    .B(_1181_),
    .X(_1339_));
 sky130_fd_sc_hd__xnor2_1 _6329_ (.A(_1239_),
    .B(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__or2_1 _6330_ (.A(_1338_),
    .B(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__nand2_1 _6331_ (.A(net30),
    .B(net35),
    .Y(_1343_));
 sky130_fd_sc_hd__xor2_1 _6332_ (.A(_1184_),
    .B(_1186_),
    .X(_1344_));
 sky130_fd_sc_hd__xnor2_1 _6333_ (.A(_1238_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__a21o_1 _6334_ (.A1(net30),
    .A2(net35),
    .B1(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__and3_1 _6335_ (.A(net30),
    .B(net35),
    .C(_1345_),
    .X(_1347_));
 sky130_fd_sc_hd__nand2_1 _6336_ (.A(net29),
    .B(net35),
    .Y(_1348_));
 sky130_fd_sc_hd__a21o_1 _6337_ (.A1(_1192_),
    .A2(_1193_),
    .B1(_1237_),
    .X(_1349_));
 sky130_fd_sc_hd__nand3_1 _6338_ (.A(_1192_),
    .B(_1193_),
    .C(_1237_),
    .Y(_1350_));
 sky130_fd_sc_hd__a21oi_1 _6339_ (.A1(_1349_),
    .A2(_1350_),
    .B1(_1348_),
    .Y(_1351_));
 sky130_fd_sc_hd__a21o_1 _6340_ (.A1(_1349_),
    .A2(_1350_),
    .B1(_1348_),
    .X(_1352_));
 sky130_fd_sc_hd__and3_1 _6341_ (.A(_1348_),
    .B(_1349_),
    .C(_1350_),
    .X(_1354_));
 sky130_fd_sc_hd__and2_1 _6342_ (.A(net28),
    .B(net35),
    .X(_1355_));
 sky130_fd_sc_hd__a211o_1 _6343_ (.A1(_1197_),
    .A2(_1200_),
    .B1(_1204_),
    .C1(_1236_),
    .X(_1356_));
 sky130_fd_sc_hd__o211ai_2 _6344_ (.A1(_1204_),
    .A2(_1236_),
    .B1(_1197_),
    .C1(_1200_),
    .Y(_1357_));
 sky130_fd_sc_hd__a21o_1 _6345_ (.A1(_1356_),
    .A2(_1357_),
    .B1(_1355_),
    .X(_1358_));
 sky130_fd_sc_hd__and3_1 _6346_ (.A(_1355_),
    .B(_1356_),
    .C(_1357_),
    .X(_1359_));
 sky130_fd_sc_hd__nand3_1 _6347_ (.A(_1355_),
    .B(_1356_),
    .C(_1357_),
    .Y(_1360_));
 sky130_fd_sc_hd__xor2_1 _6348_ (.A(_1201_),
    .B(_1203_),
    .X(_1361_));
 sky130_fd_sc_hd__xnor2_1 _6349_ (.A(_1235_),
    .B(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__nor2_1 _6350_ (.A(_4187_),
    .B(_0055_),
    .Y(_1363_));
 sky130_fd_sc_hd__or2_1 _6351_ (.A(_1362_),
    .B(_1363_),
    .X(_1365_));
 sky130_fd_sc_hd__nand2_1 _6352_ (.A(net26),
    .B(net35),
    .Y(_1366_));
 sky130_fd_sc_hd__xnor2_1 _6353_ (.A(_1205_),
    .B(_1207_),
    .Y(_1367_));
 sky130_fd_sc_hd__xnor2_1 _6354_ (.A(_1234_),
    .B(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__and3_1 _6355_ (.A(net26),
    .B(net35),
    .C(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__a21o_1 _6356_ (.A1(net26),
    .A2(net35),
    .B1(_1368_),
    .X(_1370_));
 sky130_fd_sc_hd__nand2_1 _6357_ (.A(net23),
    .B(net35),
    .Y(_1371_));
 sky130_fd_sc_hd__o22ai_2 _6358_ (.A1(_1213_),
    .A2(_1215_),
    .B1(_1220_),
    .B2(_1233_),
    .Y(_1372_));
 sky130_fd_sc_hd__or4_1 _6359_ (.A(_1213_),
    .B(_1215_),
    .C(_1220_),
    .D(_1233_),
    .X(_1373_));
 sky130_fd_sc_hd__a21oi_1 _6360_ (.A1(_1372_),
    .A2(_1373_),
    .B1(_1371_),
    .Y(_1374_));
 sky130_fd_sc_hd__a21o_1 _6361_ (.A1(_1372_),
    .A2(_1373_),
    .B1(_1371_),
    .X(_1376_));
 sky130_fd_sc_hd__and3_1 _6362_ (.A(_1371_),
    .B(_1372_),
    .C(_1373_),
    .X(_1377_));
 sky130_fd_sc_hd__and2_1 _6363_ (.A(net12),
    .B(net35),
    .X(_1378_));
 sky130_fd_sc_hd__o211ai_1 _6364_ (.A1(_1219_),
    .A2(_1220_),
    .B1(_1225_),
    .C1(_1230_),
    .Y(_1379_));
 sky130_fd_sc_hd__a211o_1 _6365_ (.A1(_1225_),
    .A2(_1230_),
    .B1(_1219_),
    .C1(_1220_),
    .X(_1380_));
 sky130_fd_sc_hd__a21oi_1 _6366_ (.A1(_1379_),
    .A2(_1380_),
    .B1(_1378_),
    .Y(_1381_));
 sky130_fd_sc_hd__nand3_1 _6367_ (.A(_1378_),
    .B(_1379_),
    .C(_1380_),
    .Y(_1382_));
 sky130_fd_sc_hd__and2b_1 _6368_ (.A_N(_1230_),
    .B(_1225_),
    .X(_1383_));
 sky130_fd_sc_hd__a21boi_1 _6369_ (.A1(_1225_),
    .A2(_1226_),
    .B1_N(_1229_),
    .Y(_1384_));
 sky130_fd_sc_hd__or4_1 _6370_ (.A(_4198_),
    .B(_0055_),
    .C(_1383_),
    .D(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__o21a_1 _6371_ (.A1(_1381_),
    .A2(_1385_),
    .B1(_1382_),
    .X(_1387_));
 sky130_fd_sc_hd__a21oi_1 _6372_ (.A1(_1376_),
    .A2(_1387_),
    .B1(_1377_),
    .Y(_1388_));
 sky130_fd_sc_hd__a21oi_1 _6373_ (.A1(_1370_),
    .A2(_1388_),
    .B1(_1369_),
    .Y(_1389_));
 sky130_fd_sc_hd__a221o_1 _6374_ (.A1(_1362_),
    .A2(_1363_),
    .B1(_1370_),
    .B2(_1388_),
    .C1(_1369_),
    .X(_1390_));
 sky130_fd_sc_hd__a31oi_1 _6375_ (.A1(_1358_),
    .A2(_1365_),
    .A3(_1390_),
    .B1(_1359_),
    .Y(_1391_));
 sky130_fd_sc_hd__a21oi_1 _6376_ (.A1(_1352_),
    .A2(_1391_),
    .B1(_1354_),
    .Y(_1392_));
 sky130_fd_sc_hd__a21oi_1 _6377_ (.A1(_1346_),
    .A2(_1392_),
    .B1(_1347_),
    .Y(_1393_));
 sky130_fd_sc_hd__a221o_1 _6378_ (.A1(_1338_),
    .A2(_1340_),
    .B1(_1346_),
    .B2(_1392_),
    .C1(_1347_),
    .X(_1394_));
 sky130_fd_sc_hd__and2_1 _6379_ (.A(_1341_),
    .B(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__o211a_1 _6380_ (.A1(_1333_),
    .A2(_1335_),
    .B1(_1341_),
    .C1(_1394_),
    .X(_1396_));
 sky130_fd_sc_hd__a22o_1 _6381_ (.A1(_1333_),
    .A2(_1335_),
    .B1(_1341_),
    .B2(_1394_),
    .X(_1398_));
 sky130_fd_sc_hd__a31o_1 _6382_ (.A1(_1329_),
    .A2(_1337_),
    .A3(_1398_),
    .B1(_1330_),
    .X(_1399_));
 sky130_fd_sc_hd__a21o_1 _6383_ (.A1(_1324_),
    .A2(_1399_),
    .B1(_1325_),
    .X(_1400_));
 sky130_fd_sc_hd__o21ai_1 _6384_ (.A1(_1319_),
    .A2(_1400_),
    .B1(_1318_),
    .Y(_1401_));
 sky130_fd_sc_hd__o221a_1 _6385_ (.A1(_1311_),
    .A2(_1313_),
    .B1(_1319_),
    .B2(_1400_),
    .C1(_1318_),
    .X(_1402_));
 sky130_fd_sc_hd__or4_2 _6386_ (.A(_1308_),
    .B(_1310_),
    .C(_1314_),
    .D(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__o22a_1 _6387_ (.A1(_1308_),
    .A2(_1310_),
    .B1(_1314_),
    .B2(_1402_),
    .X(_1404_));
 sky130_fd_sc_hd__o22ai_2 _6388_ (.A1(_1308_),
    .A2(_1310_),
    .B1(_1314_),
    .B2(_1402_),
    .Y(_1405_));
 sky130_fd_sc_hd__nand2_1 _6389_ (.A(net6),
    .B(net35),
    .Y(_1406_));
 sky130_fd_sc_hd__inv_2 _6390_ (.A(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__o41a_1 _6391_ (.A1(_1308_),
    .A2(_1310_),
    .A3(_1314_),
    .A4(_1402_),
    .B1(net35),
    .X(_1409_));
 sky130_fd_sc_hd__a211o_1 _6392_ (.A1(net6),
    .A2(_1409_),
    .B1(_1404_),
    .C1(_1307_),
    .X(_1410_));
 sky130_fd_sc_hd__xor2_1 _6393_ (.A(_1253_),
    .B(_1256_),
    .X(_1411_));
 sky130_fd_sc_hd__xnor2_1 _6394_ (.A(_1258_),
    .B(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__a21o_1 _6395_ (.A1(_1306_),
    .A2(_1410_),
    .B1(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__nand3_1 _6396_ (.A(_1306_),
    .B(_1410_),
    .C(_1412_),
    .Y(_1414_));
 sky130_fd_sc_hd__and2_1 _6397_ (.A(net8),
    .B(net35),
    .X(_1415_));
 sky130_fd_sc_hd__a31o_1 _6398_ (.A1(_1306_),
    .A2(_1410_),
    .A3(_1412_),
    .B1(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__a31o_1 _6399_ (.A1(_1301_),
    .A2(_1413_),
    .A3(_1416_),
    .B1(_1299_),
    .X(_1417_));
 sky130_fd_sc_hd__xor2_1 _6400_ (.A(_1136_),
    .B(_1260_),
    .X(_1418_));
 sky130_fd_sc_hd__xnor2_1 _6401_ (.A(_1262_),
    .B(_1418_),
    .Y(_1420_));
 sky130_fd_sc_hd__nor2_1 _6402_ (.A(_1417_),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__and2_1 _6403_ (.A(net10),
    .B(net35),
    .X(_1422_));
 sky130_fd_sc_hd__a21oi_1 _6404_ (.A1(_1417_),
    .A2(_1420_),
    .B1(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__o31ai_2 _6405_ (.A1(_1295_),
    .A2(_1421_),
    .A3(_1423_),
    .B1(_1294_),
    .Y(_1424_));
 sky130_fd_sc_hd__xor2_1 _6406_ (.A(_1264_),
    .B(_1267_),
    .X(_1425_));
 sky130_fd_sc_hd__xnor2_1 _6407_ (.A(_1269_),
    .B(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hd__or2_1 _6408_ (.A(_1424_),
    .B(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__nand2_1 _6409_ (.A(net13),
    .B(net35),
    .Y(_1428_));
 sky130_fd_sc_hd__a21bo_1 _6410_ (.A1(_1424_),
    .A2(_1426_),
    .B1_N(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__a31oi_2 _6411_ (.A1(_1288_),
    .A2(_1427_),
    .A3(_1429_),
    .B1(_1289_),
    .Y(_1431_));
 sky130_fd_sc_hd__or2_1 _6412_ (.A(_1282_),
    .B(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__nand2_1 _6413_ (.A(net15),
    .B(net35),
    .Y(_1433_));
 sky130_fd_sc_hd__a21o_1 _6414_ (.A1(_1282_),
    .A2(_1431_),
    .B1(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__nand2_1 _6415_ (.A(_1432_),
    .B(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__a21o_1 _6416_ (.A1(_1432_),
    .A2(_1434_),
    .B1(_1280_),
    .X(_1436_));
 sky130_fd_sc_hd__nand3_1 _6417_ (.A(_1280_),
    .B(_1432_),
    .C(_1434_),
    .Y(_1437_));
 sky130_fd_sc_hd__and3_1 _6418_ (.A(_3982_),
    .B(_1436_),
    .C(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__a21oi_1 _6419_ (.A1(_1436_),
    .A2(_1437_),
    .B1(_3982_),
    .Y(_1439_));
 sky130_fd_sc_hd__a21o_1 _6420_ (.A1(_1436_),
    .A2(_1437_),
    .B1(_3982_),
    .X(_1440_));
 sky130_fd_sc_hd__nor2_1 _6421_ (.A(_0000_),
    .B(_0066_),
    .Y(_1442_));
 sky130_fd_sc_hd__a2bb2o_1 _6422_ (.A1_N(_1286_),
    .A2_N(_1289_),
    .B1(_1427_),
    .B2(_1429_),
    .X(_1443_));
 sky130_fd_sc_hd__or4bb_1 _6423_ (.A(_1286_),
    .B(_1289_),
    .C_N(_1427_),
    .D_N(_1429_),
    .X(_1444_));
 sky130_fd_sc_hd__a21oi_1 _6424_ (.A1(_1443_),
    .A2(_1444_),
    .B1(_1442_),
    .Y(_1445_));
 sky130_fd_sc_hd__a21o_1 _6425_ (.A1(_1443_),
    .A2(_1444_),
    .B1(_1442_),
    .X(_1446_));
 sky130_fd_sc_hd__and3_1 _6426_ (.A(_1442_),
    .B(_1443_),
    .C(_1444_),
    .X(_1447_));
 sky130_fd_sc_hd__o22ai_1 _6427_ (.A1(_1293_),
    .A2(_1295_),
    .B1(_1421_),
    .B2(_1423_),
    .Y(_1448_));
 sky130_fd_sc_hd__or4_1 _6428_ (.A(_1293_),
    .B(_1295_),
    .C(_1421_),
    .D(_1423_),
    .X(_1449_));
 sky130_fd_sc_hd__and4_1 _6429_ (.A(net10),
    .B(net36),
    .C(_1448_),
    .D(_1449_),
    .X(_1450_));
 sky130_fd_sc_hd__a22oi_1 _6430_ (.A1(net10),
    .A2(net36),
    .B1(_1448_),
    .B2(_1449_),
    .Y(_1451_));
 sky130_fd_sc_hd__a22o_1 _6431_ (.A1(net10),
    .A2(net36),
    .B1(_1448_),
    .B2(_1449_),
    .X(_1453_));
 sky130_fd_sc_hd__a22o_1 _6432_ (.A1(_1300_),
    .A2(_1301_),
    .B1(_1413_),
    .B2(_1416_),
    .X(_1454_));
 sky130_fd_sc_hd__nand4_2 _6433_ (.A(_1300_),
    .B(_1301_),
    .C(_1413_),
    .D(_1416_),
    .Y(_1455_));
 sky130_fd_sc_hd__nand4_2 _6434_ (.A(net8),
    .B(net36),
    .C(_1454_),
    .D(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__a22oi_1 _6435_ (.A1(net8),
    .A2(net36),
    .B1(_1454_),
    .B2(_1455_),
    .Y(_1457_));
 sky130_fd_sc_hd__a22o_1 _6436_ (.A1(net8),
    .A2(net36),
    .B1(_1454_),
    .B2(_1455_),
    .X(_1458_));
 sky130_fd_sc_hd__nand2_1 _6437_ (.A(net6),
    .B(net36),
    .Y(_1459_));
 sky130_fd_sc_hd__o221ai_4 _6438_ (.A1(_1305_),
    .A2(_1307_),
    .B1(_1404_),
    .B2(_1407_),
    .C1(_1403_),
    .Y(_1460_));
 sky130_fd_sc_hd__a2111o_1 _6439_ (.A1(net6),
    .A2(_1409_),
    .B1(_1404_),
    .C1(_1307_),
    .D1(_1305_),
    .X(_1461_));
 sky130_fd_sc_hd__and3_1 _6440_ (.A(_1459_),
    .B(_1460_),
    .C(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__nand3_2 _6441_ (.A(_1459_),
    .B(_1460_),
    .C(_1461_),
    .Y(_1464_));
 sky130_fd_sc_hd__a21oi_1 _6442_ (.A1(_1460_),
    .A2(_1461_),
    .B1(_1459_),
    .Y(_1465_));
 sky130_fd_sc_hd__a21o_1 _6443_ (.A1(_1460_),
    .A2(_1461_),
    .B1(_1459_),
    .X(_1466_));
 sky130_fd_sc_hd__nand2_1 _6444_ (.A(net4),
    .B(net36),
    .Y(_1467_));
 sky130_fd_sc_hd__inv_2 _6445_ (.A(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__xor2_1 _6446_ (.A(_1311_),
    .B(_1313_),
    .X(_1469_));
 sky130_fd_sc_hd__xnor2_1 _6447_ (.A(_1401_),
    .B(_1469_),
    .Y(_1470_));
 sky130_fd_sc_hd__and2_1 _6448_ (.A(_1468_),
    .B(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__nand2_1 _6449_ (.A(net3),
    .B(net36),
    .Y(_1472_));
 sky130_fd_sc_hd__xor2_1 _6450_ (.A(_1315_),
    .B(_1317_),
    .X(_1473_));
 sky130_fd_sc_hd__xnor2_1 _6451_ (.A(_1400_),
    .B(_1473_),
    .Y(_1475_));
 sky130_fd_sc_hd__and3_1 _6452_ (.A(net3),
    .B(net36),
    .C(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__a21o_1 _6453_ (.A1(net3),
    .A2(net36),
    .B1(_1475_),
    .X(_1477_));
 sky130_fd_sc_hd__nand2_1 _6454_ (.A(net2),
    .B(net36),
    .Y(_1478_));
 sky130_fd_sc_hd__xor2_1 _6455_ (.A(_1321_),
    .B(_1323_),
    .X(_1479_));
 sky130_fd_sc_hd__xnor2_1 _6456_ (.A(_1399_),
    .B(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__and2b_1 _6457_ (.A_N(_1480_),
    .B(_1478_),
    .X(_1481_));
 sky130_fd_sc_hd__nand2b_1 _6458_ (.A_N(_1478_),
    .B(_1480_),
    .Y(_1482_));
 sky130_fd_sc_hd__and2_1 _6459_ (.A(net32),
    .B(net36),
    .X(_1483_));
 sky130_fd_sc_hd__a211o_1 _6460_ (.A1(_1329_),
    .A2(_1332_),
    .B1(_1336_),
    .C1(_1396_),
    .X(_1484_));
 sky130_fd_sc_hd__o211ai_2 _6461_ (.A1(_1336_),
    .A2(_1396_),
    .B1(_1329_),
    .C1(_1332_),
    .Y(_1486_));
 sky130_fd_sc_hd__a21oi_1 _6462_ (.A1(_1484_),
    .A2(_1486_),
    .B1(_1483_),
    .Y(_1487_));
 sky130_fd_sc_hd__a21o_1 _6463_ (.A1(_1484_),
    .A2(_1486_),
    .B1(_1483_),
    .X(_1488_));
 sky130_fd_sc_hd__and3_1 _6464_ (.A(_1483_),
    .B(_1484_),
    .C(_1486_),
    .X(_1489_));
 sky130_fd_sc_hd__nand2_1 _6465_ (.A(net31),
    .B(net36),
    .Y(_1490_));
 sky130_fd_sc_hd__inv_2 _6466_ (.A(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__xnor2_1 _6467_ (.A(_1333_),
    .B(_1335_),
    .Y(_1492_));
 sky130_fd_sc_hd__xnor2_1 _6468_ (.A(_1395_),
    .B(_1492_),
    .Y(_1493_));
 sky130_fd_sc_hd__or2_1 _6469_ (.A(_1491_),
    .B(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__nand2_1 _6470_ (.A(net30),
    .B(net36),
    .Y(_1495_));
 sky130_fd_sc_hd__xor2_1 _6471_ (.A(_1338_),
    .B(_1340_),
    .X(_1497_));
 sky130_fd_sc_hd__xnor2_1 _6472_ (.A(_1393_),
    .B(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__a21o_1 _6473_ (.A1(net30),
    .A2(net36),
    .B1(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__and3_1 _6474_ (.A(net30),
    .B(net36),
    .C(_1498_),
    .X(_1500_));
 sky130_fd_sc_hd__nand2_1 _6475_ (.A(net29),
    .B(net36),
    .Y(_1501_));
 sky130_fd_sc_hd__xor2_1 _6476_ (.A(_1343_),
    .B(_1345_),
    .X(_1502_));
 sky130_fd_sc_hd__xnor2_1 _6477_ (.A(_1392_),
    .B(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__and3_1 _6478_ (.A(net29),
    .B(net36),
    .C(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__nand2b_1 _6479_ (.A_N(_1503_),
    .B(_1501_),
    .Y(_1505_));
 sky130_fd_sc_hd__o21ai_1 _6480_ (.A1(_1351_),
    .A2(_1354_),
    .B1(_1391_),
    .Y(_1506_));
 sky130_fd_sc_hd__or3_1 _6481_ (.A(_1351_),
    .B(_1354_),
    .C(_1391_),
    .X(_1508_));
 sky130_fd_sc_hd__a22o_1 _6482_ (.A1(net28),
    .A2(net36),
    .B1(_1506_),
    .B2(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__nand4_1 _6483_ (.A(net28),
    .B(net36),
    .C(_1506_),
    .D(_1508_),
    .Y(_1510_));
 sky130_fd_sc_hd__a22o_1 _6484_ (.A1(_1358_),
    .A2(_1360_),
    .B1(_1365_),
    .B2(_1390_),
    .X(_1511_));
 sky130_fd_sc_hd__nand4_1 _6485_ (.A(_1358_),
    .B(_1360_),
    .C(_1365_),
    .D(_1390_),
    .Y(_1512_));
 sky130_fd_sc_hd__and4_1 _6486_ (.A(net27),
    .B(net36),
    .C(_1511_),
    .D(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__nand4_1 _6487_ (.A(net27),
    .B(net36),
    .C(_1511_),
    .D(_1512_),
    .Y(_1514_));
 sky130_fd_sc_hd__o2bb2a_1 _6488_ (.A1_N(_1511_),
    .A2_N(_1512_),
    .B1(_4187_),
    .B2(_0066_),
    .X(_1515_));
 sky130_fd_sc_hd__and2_1 _6489_ (.A(net26),
    .B(net36),
    .X(_1516_));
 sky130_fd_sc_hd__xor2_1 _6490_ (.A(_1362_),
    .B(_1363_),
    .X(_1517_));
 sky130_fd_sc_hd__xnor2_2 _6491_ (.A(_1389_),
    .B(_1517_),
    .Y(_1519_));
 sky130_fd_sc_hd__nand2_1 _6492_ (.A(_1516_),
    .B(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__nand2_1 _6493_ (.A(net23),
    .B(net36),
    .Y(_1521_));
 sky130_fd_sc_hd__xor2_1 _6494_ (.A(_1366_),
    .B(_1368_),
    .X(_1522_));
 sky130_fd_sc_hd__xnor2_1 _6495_ (.A(_1388_),
    .B(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__and3_1 _6496_ (.A(net23),
    .B(net36),
    .C(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__a21o_1 _6497_ (.A1(net23),
    .A2(net36),
    .B1(_1523_),
    .X(_1525_));
 sky130_fd_sc_hd__o21ai_1 _6498_ (.A1(_1374_),
    .A2(_1377_),
    .B1(_1387_),
    .Y(_1526_));
 sky130_fd_sc_hd__or3_1 _6499_ (.A(_1374_),
    .B(_1377_),
    .C(_1387_),
    .X(_1527_));
 sky130_fd_sc_hd__and4_1 _6500_ (.A(net12),
    .B(net36),
    .C(_1526_),
    .D(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__a22oi_2 _6501_ (.A1(net12),
    .A2(net36),
    .B1(_1526_),
    .B2(_1527_),
    .Y(_1530_));
 sky130_fd_sc_hd__nor2_1 _6502_ (.A(_1382_),
    .B(_1385_),
    .Y(_1531_));
 sky130_fd_sc_hd__nand2_1 _6503_ (.A(_1381_),
    .B(_1385_),
    .Y(_1532_));
 sky130_fd_sc_hd__o2111ai_4 _6504_ (.A1(_1387_),
    .A2(_1531_),
    .B1(_1532_),
    .C1(net36),
    .D1(net1),
    .Y(_1533_));
 sky130_fd_sc_hd__o21bai_2 _6505_ (.A1(_1530_),
    .A2(_1533_),
    .B1_N(_1528_),
    .Y(_1534_));
 sky130_fd_sc_hd__o21a_1 _6506_ (.A1(_1524_),
    .A2(_1534_),
    .B1(_1525_),
    .X(_1535_));
 sky130_fd_sc_hd__o221ai_4 _6507_ (.A1(_1516_),
    .A2(_1519_),
    .B1(_1524_),
    .B2(_1534_),
    .C1(_1525_),
    .Y(_1536_));
 sky130_fd_sc_hd__a31oi_2 _6508_ (.A1(_1514_),
    .A2(_1520_),
    .A3(_1536_),
    .B1(_1515_),
    .Y(_1537_));
 sky130_fd_sc_hd__a21bo_1 _6509_ (.A1(_1509_),
    .A2(_1537_),
    .B1_N(_1510_),
    .X(_1538_));
 sky130_fd_sc_hd__o21a_1 _6510_ (.A1(_1504_),
    .A2(_1538_),
    .B1(_1505_),
    .X(_1539_));
 sky130_fd_sc_hd__a21o_1 _6511_ (.A1(_1499_),
    .A2(_1539_),
    .B1(_1500_),
    .X(_1541_));
 sky130_fd_sc_hd__a221o_1 _6512_ (.A1(_1491_),
    .A2(_1493_),
    .B1(_1499_),
    .B2(_1539_),
    .C1(_1500_),
    .X(_1542_));
 sky130_fd_sc_hd__a31oi_2 _6513_ (.A1(_1488_),
    .A2(_1494_),
    .A3(_1542_),
    .B1(_1489_),
    .Y(_1543_));
 sky130_fd_sc_hd__o21ai_2 _6514_ (.A1(_1481_),
    .A2(_1543_),
    .B1(_1482_),
    .Y(_1544_));
 sky130_fd_sc_hd__o21ai_1 _6515_ (.A1(_1476_),
    .A2(_1544_),
    .B1(_1477_),
    .Y(_1545_));
 sky130_fd_sc_hd__o221a_1 _6516_ (.A1(_1468_),
    .A2(_1470_),
    .B1(_1476_),
    .B2(_1544_),
    .C1(_1477_),
    .X(_1546_));
 sky130_fd_sc_hd__and3_1 _6517_ (.A(_1403_),
    .B(_1405_),
    .C(_1406_),
    .X(_1547_));
 sky130_fd_sc_hd__a21oi_2 _6518_ (.A1(_1403_),
    .A2(_1405_),
    .B1(_1406_),
    .Y(_1548_));
 sky130_fd_sc_hd__or4_2 _6519_ (.A(_1471_),
    .B(_1546_),
    .C(_1547_),
    .D(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__o22a_2 _6520_ (.A1(_1471_),
    .A2(_1546_),
    .B1(_1547_),
    .B2(_1548_),
    .X(_1550_));
 sky130_fd_sc_hd__o22ai_2 _6521_ (.A1(_1471_),
    .A2(_1546_),
    .B1(_1547_),
    .B2(_1548_),
    .Y(_1552_));
 sky130_fd_sc_hd__and2_1 _6522_ (.A(net5),
    .B(net36),
    .X(_1553_));
 sky130_fd_sc_hd__nand2_1 _6523_ (.A(net5),
    .B(net36),
    .Y(_1554_));
 sky130_fd_sc_hd__o41a_1 _6524_ (.A1(_1471_),
    .A2(_1546_),
    .A3(_1547_),
    .A4(_1548_),
    .B1(net36),
    .X(_1555_));
 sky130_fd_sc_hd__a211oi_2 _6525_ (.A1(net5),
    .A2(_1555_),
    .B1(_1550_),
    .C1(_1465_),
    .Y(_1556_));
 sky130_fd_sc_hd__a21oi_1 _6526_ (.A1(_1413_),
    .A2(_1414_),
    .B1(_1415_),
    .Y(_1557_));
 sky130_fd_sc_hd__and3_1 _6527_ (.A(_1413_),
    .B(_1414_),
    .C(_1415_),
    .X(_1558_));
 sky130_fd_sc_hd__o22a_1 _6528_ (.A1(_1462_),
    .A2(_1556_),
    .B1(_1557_),
    .B2(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__o22ai_1 _6529_ (.A1(_1462_),
    .A2(_1556_),
    .B1(_1557_),
    .B2(_1558_),
    .Y(_1560_));
 sky130_fd_sc_hd__or4_1 _6530_ (.A(_1462_),
    .B(_1556_),
    .C(_1557_),
    .D(_1558_),
    .X(_1561_));
 sky130_fd_sc_hd__and2_1 _6531_ (.A(net7),
    .B(net36),
    .X(_1563_));
 sky130_fd_sc_hd__nand2_1 _6532_ (.A(net7),
    .B(net36),
    .Y(_1564_));
 sky130_fd_sc_hd__o41a_1 _6533_ (.A1(_1462_),
    .A2(_1556_),
    .A3(_1557_),
    .A4(_1558_),
    .B1(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__o31a_1 _6534_ (.A1(_1457_),
    .A2(_1559_),
    .A3(_1565_),
    .B1(_1456_),
    .X(_1566_));
 sky130_fd_sc_hd__xor2_1 _6535_ (.A(_1417_),
    .B(_1420_),
    .X(_1567_));
 sky130_fd_sc_hd__xnor2_1 _6536_ (.A(_1422_),
    .B(_1567_),
    .Y(_1568_));
 sky130_fd_sc_hd__nor2_1 _6537_ (.A(_1566_),
    .B(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__nand2_1 _6538_ (.A(net9),
    .B(net36),
    .Y(_1570_));
 sky130_fd_sc_hd__a21oi_1 _6539_ (.A1(_1566_),
    .A2(_1568_),
    .B1(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hd__o31a_1 _6540_ (.A1(_1450_),
    .A2(_1569_),
    .A3(_1571_),
    .B1(_1453_),
    .X(_1572_));
 sky130_fd_sc_hd__xor2_1 _6541_ (.A(_1424_),
    .B(_1426_),
    .X(_1574_));
 sky130_fd_sc_hd__xnor2_1 _6542_ (.A(_1428_),
    .B(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hd__or2_1 _6543_ (.A(_1572_),
    .B(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__and2_1 _6544_ (.A(net11),
    .B(net36),
    .X(_1577_));
 sky130_fd_sc_hd__a21o_1 _6545_ (.A1(_1572_),
    .A2(_1575_),
    .B1(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__a31o_1 _6546_ (.A1(_1446_),
    .A2(_1576_),
    .A3(_1578_),
    .B1(_1447_),
    .X(_1579_));
 sky130_fd_sc_hd__xor2_1 _6547_ (.A(_1282_),
    .B(_1431_),
    .X(_1580_));
 sky130_fd_sc_hd__xnor2_2 _6548_ (.A(_1433_),
    .B(_1580_),
    .Y(_1581_));
 sky130_fd_sc_hd__nor2_1 _6549_ (.A(_1579_),
    .B(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__and2_1 _6550_ (.A(net14),
    .B(net36),
    .X(_1583_));
 sky130_fd_sc_hd__a21oi_1 _6551_ (.A1(_1579_),
    .A2(_1581_),
    .B1(_1583_),
    .Y(_1585_));
 sky130_fd_sc_hd__o31a_1 _6552_ (.A1(_1438_),
    .A2(_1582_),
    .A3(_1585_),
    .B1(_1440_),
    .X(_1586_));
 sky130_fd_sc_hd__a21boi_2 _6553_ (.A1(_1278_),
    .A2(_1435_),
    .B1_N(_1279_),
    .Y(_1587_));
 sky130_fd_sc_hd__a21oi_2 _6554_ (.A1(_1586_),
    .A2(_1587_),
    .B1(_3981_),
    .Y(_1588_));
 sky130_fd_sc_hd__a21o_1 _6555_ (.A1(net37),
    .A2(_1716_),
    .B1(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__a21bo_1 _6556_ (.A1(net37),
    .A2(_1588_),
    .B1_N(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__xor2_1 _6557_ (.A(_1586_),
    .B(_1587_),
    .X(_1591_));
 sky130_fd_sc_hd__xnor2_2 _6558_ (.A(_3981_),
    .B(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__and2_1 _6559_ (.A(net14),
    .B(net37),
    .X(_1593_));
 sky130_fd_sc_hd__o22ai_1 _6560_ (.A1(_1438_),
    .A2(_1439_),
    .B1(_1582_),
    .B2(_1585_),
    .Y(_1594_));
 sky130_fd_sc_hd__or4_1 _6561_ (.A(_1438_),
    .B(_1439_),
    .C(_1582_),
    .D(_1585_),
    .X(_1596_));
 sky130_fd_sc_hd__and3_1 _6562_ (.A(_1593_),
    .B(_1594_),
    .C(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__a21oi_1 _6563_ (.A1(_1594_),
    .A2(_1596_),
    .B1(_1593_),
    .Y(_1598_));
 sky130_fd_sc_hd__a21o_1 _6564_ (.A1(_1594_),
    .A2(_1596_),
    .B1(_1593_),
    .X(_1599_));
 sky130_fd_sc_hd__nand2_1 _6565_ (.A(net11),
    .B(net37),
    .Y(_1600_));
 sky130_fd_sc_hd__o211ai_2 _6566_ (.A1(_1445_),
    .A2(_1447_),
    .B1(_1576_),
    .C1(_1578_),
    .Y(_1601_));
 sky130_fd_sc_hd__a211o_1 _6567_ (.A1(_1576_),
    .A2(_1578_),
    .B1(_1445_),
    .C1(_1447_),
    .X(_1602_));
 sky130_fd_sc_hd__nand3_1 _6568_ (.A(_1600_),
    .B(_1601_),
    .C(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__a21oi_1 _6569_ (.A1(_1601_),
    .A2(_1602_),
    .B1(_1600_),
    .Y(_1604_));
 sky130_fd_sc_hd__a21o_1 _6570_ (.A1(_1601_),
    .A2(_1602_),
    .B1(_1600_),
    .X(_1605_));
 sky130_fd_sc_hd__nand2_1 _6571_ (.A(net9),
    .B(net37),
    .Y(_1607_));
 sky130_fd_sc_hd__o22ai_1 _6572_ (.A1(_1450_),
    .A2(_1451_),
    .B1(_1569_),
    .B2(_1571_),
    .Y(_1608_));
 sky130_fd_sc_hd__or4_1 _6573_ (.A(_1450_),
    .B(_1451_),
    .C(_1569_),
    .D(_1571_),
    .X(_1609_));
 sky130_fd_sc_hd__and3_1 _6574_ (.A(_1607_),
    .B(_1608_),
    .C(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__nand3_1 _6575_ (.A(_1607_),
    .B(_1608_),
    .C(_1609_),
    .Y(_1611_));
 sky130_fd_sc_hd__a21oi_1 _6576_ (.A1(_1608_),
    .A2(_1609_),
    .B1(_1607_),
    .Y(_1612_));
 sky130_fd_sc_hd__nand2_1 _6577_ (.A(net7),
    .B(net37),
    .Y(_1613_));
 sky130_fd_sc_hd__a211o_1 _6578_ (.A1(_1456_),
    .A2(_1458_),
    .B1(_1559_),
    .C1(_1565_),
    .X(_1614_));
 sky130_fd_sc_hd__o211ai_2 _6579_ (.A1(_1559_),
    .A2(_1565_),
    .B1(_1456_),
    .C1(_1458_),
    .Y(_1615_));
 sky130_fd_sc_hd__a21oi_1 _6580_ (.A1(_1614_),
    .A2(_1615_),
    .B1(_1613_),
    .Y(_1616_));
 sky130_fd_sc_hd__and3_1 _6581_ (.A(_1613_),
    .B(_1614_),
    .C(_1615_),
    .X(_1618_));
 sky130_fd_sc_hd__nand3_1 _6582_ (.A(_1613_),
    .B(_1614_),
    .C(_1615_),
    .Y(_1619_));
 sky130_fd_sc_hd__and2_1 _6583_ (.A(net5),
    .B(net37),
    .X(_1620_));
 sky130_fd_sc_hd__a221o_1 _6584_ (.A1(_1464_),
    .A2(_1466_),
    .B1(_1555_),
    .B2(net5),
    .C1(_1550_),
    .X(_1621_));
 sky130_fd_sc_hd__o2111ai_4 _6585_ (.A1(_1550_),
    .A2(_1553_),
    .B1(_1464_),
    .C1(_1466_),
    .D1(_1549_),
    .Y(_1622_));
 sky130_fd_sc_hd__a21oi_4 _6586_ (.A1(_1621_),
    .A2(_1622_),
    .B1(_1620_),
    .Y(_1623_));
 sky130_fd_sc_hd__and3_1 _6587_ (.A(_1620_),
    .B(_1621_),
    .C(_1622_),
    .X(_1624_));
 sky130_fd_sc_hd__nand2_1 _6588_ (.A(net3),
    .B(net37),
    .Y(_1625_));
 sky130_fd_sc_hd__inv_2 _6589_ (.A(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__xnor2_1 _6590_ (.A(_1467_),
    .B(_1470_),
    .Y(_1627_));
 sky130_fd_sc_hd__xnor2_1 _6591_ (.A(_1545_),
    .B(_1627_),
    .Y(_1629_));
 sky130_fd_sc_hd__or2_1 _6592_ (.A(_1626_),
    .B(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__nand2_1 _6593_ (.A(net2),
    .B(net37),
    .Y(_1631_));
 sky130_fd_sc_hd__xor2_1 _6594_ (.A(_1472_),
    .B(_1475_),
    .X(_1632_));
 sky130_fd_sc_hd__xnor2_1 _6595_ (.A(_1544_),
    .B(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__a21o_1 _6596_ (.A1(net2),
    .A2(net37),
    .B1(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__and3_1 _6597_ (.A(net2),
    .B(net37),
    .C(_1633_),
    .X(_1635_));
 sky130_fd_sc_hd__nand2_1 _6598_ (.A(net32),
    .B(net37),
    .Y(_1636_));
 sky130_fd_sc_hd__xnor2_1 _6599_ (.A(_1478_),
    .B(_1480_),
    .Y(_1637_));
 sky130_fd_sc_hd__xnor2_1 _6600_ (.A(_1543_),
    .B(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__and2b_1 _6601_ (.A_N(_1638_),
    .B(_1636_),
    .X(_1640_));
 sky130_fd_sc_hd__nand2b_1 _6602_ (.A_N(_1636_),
    .B(_1638_),
    .Y(_1641_));
 sky130_fd_sc_hd__nand2_1 _6603_ (.A(net31),
    .B(net37),
    .Y(_1642_));
 sky130_fd_sc_hd__a211o_1 _6604_ (.A1(_1494_),
    .A2(_1542_),
    .B1(_1487_),
    .C1(_1489_),
    .X(_1643_));
 sky130_fd_sc_hd__o211ai_2 _6605_ (.A1(_1487_),
    .A2(_1489_),
    .B1(_1494_),
    .C1(_1542_),
    .Y(_1644_));
 sky130_fd_sc_hd__and3_1 _6606_ (.A(_1642_),
    .B(_1643_),
    .C(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__a21oi_1 _6607_ (.A1(_1643_),
    .A2(_1644_),
    .B1(_1642_),
    .Y(_1646_));
 sky130_fd_sc_hd__a21o_1 _6608_ (.A1(_1643_),
    .A2(_1644_),
    .B1(_1642_),
    .X(_1647_));
 sky130_fd_sc_hd__nand2_1 _6609_ (.A(net30),
    .B(net37),
    .Y(_1648_));
 sky130_fd_sc_hd__xnor2_1 _6610_ (.A(_1490_),
    .B(_1493_),
    .Y(_1649_));
 sky130_fd_sc_hd__xnor2_1 _6611_ (.A(_1541_),
    .B(_1649_),
    .Y(_1651_));
 sky130_fd_sc_hd__and2_1 _6612_ (.A(_1648_),
    .B(_1651_),
    .X(_1652_));
 sky130_fd_sc_hd__nand2_1 _6613_ (.A(net29),
    .B(net37),
    .Y(_1653_));
 sky130_fd_sc_hd__xnor2_1 _6614_ (.A(_1495_),
    .B(_1498_),
    .Y(_1654_));
 sky130_fd_sc_hd__xnor2_1 _6615_ (.A(_1539_),
    .B(_1654_),
    .Y(_1655_));
 sky130_fd_sc_hd__and2_1 _6616_ (.A(_1653_),
    .B(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__nand2_1 _6617_ (.A(net28),
    .B(net37),
    .Y(_1657_));
 sky130_fd_sc_hd__inv_2 _6618_ (.A(_1657_),
    .Y(_1658_));
 sky130_fd_sc_hd__xor2_1 _6619_ (.A(_1501_),
    .B(_1503_),
    .X(_1659_));
 sky130_fd_sc_hd__xnor2_2 _6620_ (.A(_1538_),
    .B(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__nand2_1 _6621_ (.A(_1658_),
    .B(_1660_),
    .Y(_1662_));
 sky130_fd_sc_hd__a21o_1 _6622_ (.A1(_1509_),
    .A2(_1510_),
    .B1(_1537_),
    .X(_1663_));
 sky130_fd_sc_hd__nand3_1 _6623_ (.A(_1509_),
    .B(_1510_),
    .C(_1537_),
    .Y(_1664_));
 sky130_fd_sc_hd__and4_1 _6624_ (.A(net27),
    .B(net37),
    .C(_1663_),
    .D(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__o2bb2a_1 _6625_ (.A1_N(_1663_),
    .A2_N(_1664_),
    .B1(_4187_),
    .B2(_0077_),
    .X(_1666_));
 sky130_fd_sc_hd__a22o_1 _6626_ (.A1(net27),
    .A2(net37),
    .B1(_1663_),
    .B2(_1664_),
    .X(_1667_));
 sky130_fd_sc_hd__o211ai_2 _6627_ (.A1(_1513_),
    .A2(_1515_),
    .B1(_1520_),
    .C1(_1536_),
    .Y(_1668_));
 sky130_fd_sc_hd__a211o_1 _6628_ (.A1(_1520_),
    .A2(_1536_),
    .B1(_1513_),
    .C1(_1515_),
    .X(_1669_));
 sky130_fd_sc_hd__and2_1 _6629_ (.A(net26),
    .B(net37),
    .X(_1670_));
 sky130_fd_sc_hd__a21oi_1 _6630_ (.A1(_1668_),
    .A2(_1669_),
    .B1(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__a21o_1 _6631_ (.A1(_1668_),
    .A2(_1669_),
    .B1(_1670_),
    .X(_1673_));
 sky130_fd_sc_hd__and3_1 _6632_ (.A(_1668_),
    .B(_1669_),
    .C(_1670_),
    .X(_1674_));
 sky130_fd_sc_hd__nand2_1 _6633_ (.A(net23),
    .B(net37),
    .Y(_1675_));
 sky130_fd_sc_hd__xnor2_1 _6634_ (.A(_1516_),
    .B(_1519_),
    .Y(_1676_));
 sky130_fd_sc_hd__xnor2_1 _6635_ (.A(_1535_),
    .B(_1676_),
    .Y(_1677_));
 sky130_fd_sc_hd__nand2b_1 _6636_ (.A_N(_1677_),
    .B(_1675_),
    .Y(_1678_));
 sky130_fd_sc_hd__nand2_1 _6637_ (.A(net12),
    .B(net37),
    .Y(_1679_));
 sky130_fd_sc_hd__xnor2_1 _6638_ (.A(_1521_),
    .B(_1523_),
    .Y(_1680_));
 sky130_fd_sc_hd__xnor2_1 _6639_ (.A(_1534_),
    .B(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__nand2_1 _6640_ (.A(_1679_),
    .B(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__nor2_1 _6641_ (.A(_1679_),
    .B(_1681_),
    .Y(_1684_));
 sky130_fd_sc_hd__or2_1 _6642_ (.A(_1528_),
    .B(_1530_),
    .X(_1685_));
 sky130_fd_sc_hd__xnor2_1 _6643_ (.A(_1533_),
    .B(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__nor3_1 _6644_ (.A(_4198_),
    .B(_0077_),
    .C(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__a2111oi_1 _6645_ (.A1(_1679_),
    .A2(_1681_),
    .B1(_1686_),
    .C1(_0077_),
    .D1(_4198_),
    .Y(_1688_));
 sky130_fd_sc_hd__nor2_1 _6646_ (.A(_1684_),
    .B(_1688_),
    .Y(_1689_));
 sky130_fd_sc_hd__a311o_1 _6647_ (.A1(net23),
    .A2(net37),
    .A3(_1677_),
    .B1(_1684_),
    .C1(_1688_),
    .X(_1690_));
 sky130_fd_sc_hd__a31o_1 _6648_ (.A1(_1673_),
    .A2(_1678_),
    .A3(_1690_),
    .B1(_1674_),
    .X(_1691_));
 sky130_fd_sc_hd__o21ai_1 _6649_ (.A1(_1665_),
    .A2(_1691_),
    .B1(_1667_),
    .Y(_1692_));
 sky130_fd_sc_hd__o221ai_2 _6650_ (.A1(_1658_),
    .A2(_1660_),
    .B1(_1665_),
    .B2(_1691_),
    .C1(_1667_),
    .Y(_1693_));
 sky130_fd_sc_hd__nand2_1 _6651_ (.A(_1662_),
    .B(_1693_),
    .Y(_1695_));
 sky130_fd_sc_hd__o211a_1 _6652_ (.A1(_1653_),
    .A2(_1655_),
    .B1(_1662_),
    .C1(_1693_),
    .X(_1696_));
 sky130_fd_sc_hd__nor2_1 _6653_ (.A(_1656_),
    .B(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__o22a_1 _6654_ (.A1(_1648_),
    .A2(_1651_),
    .B1(_1656_),
    .B2(_1696_),
    .X(_1698_));
 sky130_fd_sc_hd__o31a_1 _6655_ (.A1(_1645_),
    .A2(_1652_),
    .A3(_1698_),
    .B1(_1647_),
    .X(_1699_));
 sky130_fd_sc_hd__o21ai_2 _6656_ (.A1(_1640_),
    .A2(_1699_),
    .B1(_1641_),
    .Y(_1700_));
 sky130_fd_sc_hd__a21oi_1 _6657_ (.A1(_1634_),
    .A2(_1700_),
    .B1(_1635_),
    .Y(_1701_));
 sky130_fd_sc_hd__a221o_1 _6658_ (.A1(_1626_),
    .A2(_1629_),
    .B1(_1634_),
    .B2(_1700_),
    .C1(_1635_),
    .X(_1702_));
 sky130_fd_sc_hd__and3_1 _6659_ (.A(_1549_),
    .B(_1552_),
    .C(_1554_),
    .X(_1703_));
 sky130_fd_sc_hd__a21oi_1 _6660_ (.A1(_1549_),
    .A2(_1552_),
    .B1(_1554_),
    .Y(_1704_));
 sky130_fd_sc_hd__a21o_1 _6661_ (.A1(_1549_),
    .A2(_1552_),
    .B1(_1553_),
    .X(_1706_));
 sky130_fd_sc_hd__nand4_1 _6662_ (.A(net5),
    .B(net36),
    .C(_1549_),
    .D(_1552_),
    .Y(_1707_));
 sky130_fd_sc_hd__a211o_1 _6663_ (.A1(_1630_),
    .A2(_1702_),
    .B1(_1703_),
    .C1(_1704_),
    .X(_1708_));
 sky130_fd_sc_hd__o211ai_1 _6664_ (.A1(_1703_),
    .A2(_1704_),
    .B1(_1630_),
    .C1(_1702_),
    .Y(_1709_));
 sky130_fd_sc_hd__nand2_1 _6665_ (.A(net4),
    .B(net37),
    .Y(_1710_));
 sky130_fd_sc_hd__inv_2 _6666_ (.A(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__a41o_1 _6667_ (.A1(_1630_),
    .A2(_1702_),
    .A3(_1706_),
    .A4(_1707_),
    .B1(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__a21oi_2 _6668_ (.A1(_1708_),
    .A2(_1712_),
    .B1(_1624_),
    .Y(_1713_));
 sky130_fd_sc_hd__a21oi_2 _6669_ (.A1(_1560_),
    .A2(_1561_),
    .B1(_1563_),
    .Y(_1714_));
 sky130_fd_sc_hd__and3_1 _6670_ (.A(_1560_),
    .B(_1561_),
    .C(_1563_),
    .X(_1715_));
 sky130_fd_sc_hd__o22ai_4 _6671_ (.A1(_1623_),
    .A2(_1713_),
    .B1(_1714_),
    .B2(_1715_),
    .Y(_1717_));
 sky130_fd_sc_hd__or4_1 _6672_ (.A(_1623_),
    .B(_1713_),
    .C(_1714_),
    .D(_1715_),
    .X(_1718_));
 sky130_fd_sc_hd__and2_1 _6673_ (.A(net6),
    .B(net37),
    .X(_1719_));
 sky130_fd_sc_hd__nand2_1 _6674_ (.A(net6),
    .B(net37),
    .Y(_1720_));
 sky130_fd_sc_hd__o41ai_2 _6675_ (.A1(_1623_),
    .A2(_1713_),
    .A3(_1714_),
    .A4(_1715_),
    .B1(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__a31o_1 _6676_ (.A1(_1619_),
    .A2(_1717_),
    .A3(_1721_),
    .B1(_1616_),
    .X(_1722_));
 sky130_fd_sc_hd__xor2_1 _6677_ (.A(_1566_),
    .B(_1568_),
    .X(_1723_));
 sky130_fd_sc_hd__xnor2_1 _6678_ (.A(_1570_),
    .B(_1723_),
    .Y(_1724_));
 sky130_fd_sc_hd__or2_1 _6679_ (.A(_1722_),
    .B(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__nand2_1 _6680_ (.A(net8),
    .B(net37),
    .Y(_1726_));
 sky130_fd_sc_hd__a21bo_1 _6681_ (.A1(_1722_),
    .A2(_1724_),
    .B1_N(_1726_),
    .X(_1728_));
 sky130_fd_sc_hd__a31o_1 _6682_ (.A1(_1611_),
    .A2(_1725_),
    .A3(_1728_),
    .B1(_1612_),
    .X(_1729_));
 sky130_fd_sc_hd__xnor2_1 _6683_ (.A(_1572_),
    .B(_1575_),
    .Y(_1730_));
 sky130_fd_sc_hd__xnor2_1 _6684_ (.A(_1577_),
    .B(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__or2_1 _6685_ (.A(_1729_),
    .B(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__nand2_1 _6686_ (.A(net10),
    .B(net37),
    .Y(_1733_));
 sky130_fd_sc_hd__a21bo_1 _6687_ (.A1(_1729_),
    .A2(_1731_),
    .B1_N(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__a31o_1 _6688_ (.A1(_1603_),
    .A2(_1732_),
    .A3(_1734_),
    .B1(_1604_),
    .X(_1735_));
 sky130_fd_sc_hd__xnor2_1 _6689_ (.A(_1579_),
    .B(_1581_),
    .Y(_1736_));
 sky130_fd_sc_hd__xnor2_2 _6690_ (.A(_1583_),
    .B(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__or2_1 _6691_ (.A(_1735_),
    .B(_1737_),
    .X(_1739_));
 sky130_fd_sc_hd__nand2_1 _6692_ (.A(net13),
    .B(net37),
    .Y(_1740_));
 sky130_fd_sc_hd__a21bo_1 _6693_ (.A1(_1735_),
    .A2(_1737_),
    .B1_N(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__a31o_1 _6694_ (.A1(_1599_),
    .A2(_1739_),
    .A3(_1741_),
    .B1(_1597_),
    .X(_1742_));
 sky130_fd_sc_hd__or2_1 _6695_ (.A(_1592_),
    .B(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__nand2_1 _6696_ (.A(net15),
    .B(net37),
    .Y(_1744_));
 sky130_fd_sc_hd__a21bo_1 _6697_ (.A1(_1592_),
    .A2(_1742_),
    .B1_N(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__nand3_1 _6698_ (.A(_1590_),
    .B(_1743_),
    .C(_1745_),
    .Y(_1746_));
 sky130_fd_sc_hd__a21o_1 _6699_ (.A1(_1743_),
    .A2(_1745_),
    .B1(_1590_),
    .X(_1747_));
 sky130_fd_sc_hd__and3_1 _6700_ (.A(_3980_),
    .B(_1746_),
    .C(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__a21oi_1 _6701_ (.A1(_1746_),
    .A2(_1747_),
    .B1(_3980_),
    .Y(_1750_));
 sky130_fd_sc_hd__a21o_1 _6702_ (.A1(_1746_),
    .A2(_1747_),
    .B1(_3980_),
    .X(_1751_));
 sky130_fd_sc_hd__nand2_1 _6703_ (.A(net13),
    .B(net38),
    .Y(_1752_));
 sky130_fd_sc_hd__o211ai_2 _6704_ (.A1(_1597_),
    .A2(_1598_),
    .B1(_1739_),
    .C1(_1741_),
    .Y(_1753_));
 sky130_fd_sc_hd__a211o_1 _6705_ (.A1(_1739_),
    .A2(_1741_),
    .B1(_1597_),
    .C1(_1598_),
    .X(_1754_));
 sky130_fd_sc_hd__a21oi_1 _6706_ (.A1(_1753_),
    .A2(_1754_),
    .B1(_1752_),
    .Y(_1755_));
 sky130_fd_sc_hd__a21o_1 _6707_ (.A1(_1753_),
    .A2(_1754_),
    .B1(_1752_),
    .X(_1756_));
 sky130_fd_sc_hd__nand3_1 _6708_ (.A(_1752_),
    .B(_1753_),
    .C(_1754_),
    .Y(_1757_));
 sky130_fd_sc_hd__and2_1 _6709_ (.A(net10),
    .B(net38),
    .X(_1758_));
 sky130_fd_sc_hd__a22o_1 _6710_ (.A1(_1603_),
    .A2(_1605_),
    .B1(_1732_),
    .B2(_1734_),
    .X(_1759_));
 sky130_fd_sc_hd__nand4_2 _6711_ (.A(_1603_),
    .B(_1605_),
    .C(_1732_),
    .D(_1734_),
    .Y(_1761_));
 sky130_fd_sc_hd__a21oi_2 _6712_ (.A1(_1759_),
    .A2(_1761_),
    .B1(_1758_),
    .Y(_1762_));
 sky130_fd_sc_hd__and3_1 _6713_ (.A(_1758_),
    .B(_1759_),
    .C(_1761_),
    .X(_1763_));
 sky130_fd_sc_hd__nand3_1 _6714_ (.A(_1758_),
    .B(_1759_),
    .C(_1761_),
    .Y(_1764_));
 sky130_fd_sc_hd__and2_1 _6715_ (.A(net8),
    .B(net38),
    .X(_1765_));
 sky130_fd_sc_hd__a2bb2o_1 _6716_ (.A1_N(_1610_),
    .A2_N(_1612_),
    .B1(_1725_),
    .B2(_1728_),
    .X(_1766_));
 sky130_fd_sc_hd__or4bb_1 _6717_ (.A(_1610_),
    .B(_1612_),
    .C_N(_1725_),
    .D_N(_1728_),
    .X(_1767_));
 sky130_fd_sc_hd__a21o_1 _6718_ (.A1(_1766_),
    .A2(_1767_),
    .B1(_1765_),
    .X(_1768_));
 sky130_fd_sc_hd__and3_1 _6719_ (.A(_1765_),
    .B(_1766_),
    .C(_1767_),
    .X(_1769_));
 sky130_fd_sc_hd__nand3_1 _6720_ (.A(_1765_),
    .B(_1766_),
    .C(_1767_),
    .Y(_1770_));
 sky130_fd_sc_hd__nand2_1 _6721_ (.A(net6),
    .B(net38),
    .Y(_1772_));
 sky130_fd_sc_hd__o211ai_2 _6722_ (.A1(_1616_),
    .A2(_1618_),
    .B1(_1717_),
    .C1(_1721_),
    .Y(_1773_));
 sky130_fd_sc_hd__a211o_1 _6723_ (.A1(_1717_),
    .A2(_1721_),
    .B1(_1616_),
    .C1(_1618_),
    .X(_1774_));
 sky130_fd_sc_hd__and3_1 _6724_ (.A(_1772_),
    .B(_1773_),
    .C(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__nand3_1 _6725_ (.A(_1772_),
    .B(_1773_),
    .C(_1774_),
    .Y(_1776_));
 sky130_fd_sc_hd__a21oi_1 _6726_ (.A1(_1773_),
    .A2(_1774_),
    .B1(_1772_),
    .Y(_1777_));
 sky130_fd_sc_hd__a21o_1 _6727_ (.A1(_1717_),
    .A2(_1718_),
    .B1(_1719_),
    .X(_1778_));
 sky130_fd_sc_hd__nand3_1 _6728_ (.A(_1717_),
    .B(_1718_),
    .C(_1719_),
    .Y(_1779_));
 sky130_fd_sc_hd__nand2_1 _6729_ (.A(net4),
    .B(net38),
    .Y(_1780_));
 sky130_fd_sc_hd__o211ai_2 _6730_ (.A1(_1623_),
    .A2(_1624_),
    .B1(_1708_),
    .C1(_1712_),
    .Y(_1781_));
 sky130_fd_sc_hd__a211o_1 _6731_ (.A1(_1708_),
    .A2(_1712_),
    .B1(_1623_),
    .C1(_1624_),
    .X(_1783_));
 sky130_fd_sc_hd__and3_1 _6732_ (.A(_1780_),
    .B(_1781_),
    .C(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__nand3_1 _6733_ (.A(_1780_),
    .B(_1781_),
    .C(_1783_),
    .Y(_1785_));
 sky130_fd_sc_hd__a21oi_1 _6734_ (.A1(_1781_),
    .A2(_1783_),
    .B1(_1780_),
    .Y(_1786_));
 sky130_fd_sc_hd__nand2_1 _6735_ (.A(net2),
    .B(net38),
    .Y(_1787_));
 sky130_fd_sc_hd__inv_2 _6736_ (.A(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hd__xnor2_1 _6737_ (.A(_1625_),
    .B(_1629_),
    .Y(_1789_));
 sky130_fd_sc_hd__xnor2_1 _6738_ (.A(_1701_),
    .B(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__and2_1 _6739_ (.A(_1788_),
    .B(_1790_),
    .X(_1791_));
 sky130_fd_sc_hd__nand2_1 _6740_ (.A(net32),
    .B(net38),
    .Y(_1792_));
 sky130_fd_sc_hd__xnor2_1 _6741_ (.A(_1631_),
    .B(_1633_),
    .Y(_1794_));
 sky130_fd_sc_hd__xnor2_1 _6742_ (.A(_1700_),
    .B(_1794_),
    .Y(_1795_));
 sky130_fd_sc_hd__or2_1 _6743_ (.A(_1792_),
    .B(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__nand2_1 _6744_ (.A(net31),
    .B(net38),
    .Y(_1797_));
 sky130_fd_sc_hd__xnor2_1 _6745_ (.A(_1636_),
    .B(_1638_),
    .Y(_1798_));
 sky130_fd_sc_hd__xnor2_1 _6746_ (.A(_1699_),
    .B(_1798_),
    .Y(_1799_));
 sky130_fd_sc_hd__nand2b_1 _6747_ (.A_N(_1797_),
    .B(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__a21oi_1 _6748_ (.A1(net31),
    .A2(net38),
    .B1(_1799_),
    .Y(_1801_));
 sky130_fd_sc_hd__and2_1 _6749_ (.A(net30),
    .B(net38),
    .X(_1802_));
 sky130_fd_sc_hd__o22ai_2 _6750_ (.A1(_1645_),
    .A2(_1646_),
    .B1(_1652_),
    .B2(_1698_),
    .Y(_1803_));
 sky130_fd_sc_hd__or4_1 _6751_ (.A(_1645_),
    .B(_1646_),
    .C(_1652_),
    .D(_1698_),
    .X(_1805_));
 sky130_fd_sc_hd__and3_1 _6752_ (.A(_1802_),
    .B(_1803_),
    .C(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__nand3_1 _6753_ (.A(_1802_),
    .B(_1803_),
    .C(_1805_),
    .Y(_1807_));
 sky130_fd_sc_hd__a21oi_1 _6754_ (.A1(_1803_),
    .A2(_1805_),
    .B1(_1802_),
    .Y(_1808_));
 sky130_fd_sc_hd__and2_1 _6755_ (.A(net29),
    .B(net38),
    .X(_1809_));
 sky130_fd_sc_hd__xnor2_1 _6756_ (.A(_1648_),
    .B(_1651_),
    .Y(_1810_));
 sky130_fd_sc_hd__xnor2_2 _6757_ (.A(_1697_),
    .B(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__nand2_1 _6758_ (.A(_1809_),
    .B(_1811_),
    .Y(_1812_));
 sky130_fd_sc_hd__nand2_1 _6759_ (.A(net28),
    .B(net38),
    .Y(_1813_));
 sky130_fd_sc_hd__inv_2 _6760_ (.A(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hd__xnor2_1 _6761_ (.A(_1653_),
    .B(_1655_),
    .Y(_1816_));
 sky130_fd_sc_hd__xnor2_1 _6762_ (.A(_1695_),
    .B(_1816_),
    .Y(_1817_));
 sky130_fd_sc_hd__and2_1 _6763_ (.A(_1814_),
    .B(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__nand2_1 _6764_ (.A(net27),
    .B(net38),
    .Y(_1819_));
 sky130_fd_sc_hd__xnor2_1 _6765_ (.A(_1657_),
    .B(_1660_),
    .Y(_1820_));
 sky130_fd_sc_hd__xnor2_1 _6766_ (.A(_1692_),
    .B(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__and3_1 _6767_ (.A(net27),
    .B(net38),
    .C(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__nand2b_1 _6768_ (.A_N(_1821_),
    .B(_1819_),
    .Y(_1823_));
 sky130_fd_sc_hd__o21bai_1 _6769_ (.A1(_1665_),
    .A2(_1666_),
    .B1_N(_1691_),
    .Y(_1824_));
 sky130_fd_sc_hd__or3b_1 _6770_ (.A(_1665_),
    .B(_1666_),
    .C_N(_1691_),
    .X(_1825_));
 sky130_fd_sc_hd__a22o_1 _6771_ (.A1(net26),
    .A2(net38),
    .B1(_1824_),
    .B2(_1825_),
    .X(_1827_));
 sky130_fd_sc_hd__nand4_1 _6772_ (.A(net26),
    .B(net38),
    .C(_1824_),
    .D(_1825_),
    .Y(_1828_));
 sky130_fd_sc_hd__nand2_1 _6773_ (.A(net23),
    .B(net38),
    .Y(_1829_));
 sky130_fd_sc_hd__o211ai_2 _6774_ (.A1(_1671_),
    .A2(_1674_),
    .B1(_1678_),
    .C1(_1690_),
    .Y(_1830_));
 sky130_fd_sc_hd__a211o_1 _6775_ (.A1(_1678_),
    .A2(_1690_),
    .B1(_1671_),
    .C1(_1674_),
    .X(_1831_));
 sky130_fd_sc_hd__a21oi_1 _6776_ (.A1(_1830_),
    .A2(_1831_),
    .B1(_1829_),
    .Y(_1832_));
 sky130_fd_sc_hd__a21o_1 _6777_ (.A1(_1830_),
    .A2(_1831_),
    .B1(_1829_),
    .X(_1833_));
 sky130_fd_sc_hd__and3_1 _6778_ (.A(_1829_),
    .B(_1830_),
    .C(_1831_),
    .X(_1834_));
 sky130_fd_sc_hd__and2_1 _6779_ (.A(net12),
    .B(net38),
    .X(_1835_));
 sky130_fd_sc_hd__xnor2_1 _6780_ (.A(_1675_),
    .B(_1677_),
    .Y(_1836_));
 sky130_fd_sc_hd__xnor2_1 _6781_ (.A(_1689_),
    .B(_1836_),
    .Y(_1838_));
 sky130_fd_sc_hd__nand2_1 _6782_ (.A(_1835_),
    .B(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__and2_1 _6783_ (.A(_1684_),
    .B(_1687_),
    .X(_1840_));
 sky130_fd_sc_hd__or2_1 _6784_ (.A(_1682_),
    .B(_1687_),
    .X(_1841_));
 sky130_fd_sc_hd__o2111ai_2 _6785_ (.A1(_1689_),
    .A2(_1840_),
    .B1(_1841_),
    .C1(net38),
    .D1(net1),
    .Y(_1842_));
 sky130_fd_sc_hd__o21bai_1 _6786_ (.A1(_1835_),
    .A2(_1838_),
    .B1_N(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__a31oi_2 _6787_ (.A1(_1833_),
    .A2(_1839_),
    .A3(_1843_),
    .B1(_1834_),
    .Y(_1844_));
 sky130_fd_sc_hd__a21bo_1 _6788_ (.A1(_1827_),
    .A2(_1844_),
    .B1_N(_1828_),
    .X(_1845_));
 sky130_fd_sc_hd__o21ai_1 _6789_ (.A1(_1822_),
    .A2(_1845_),
    .B1(_1823_),
    .Y(_1846_));
 sky130_fd_sc_hd__o221a_1 _6790_ (.A1(_1814_),
    .A2(_1817_),
    .B1(_1822_),
    .B2(_1845_),
    .C1(_1823_),
    .X(_1847_));
 sky130_fd_sc_hd__or2_1 _6791_ (.A(_1818_),
    .B(_1847_),
    .X(_1849_));
 sky130_fd_sc_hd__o22ai_2 _6792_ (.A1(_1809_),
    .A2(_1811_),
    .B1(_1818_),
    .B2(_1847_),
    .Y(_1850_));
 sky130_fd_sc_hd__a31o_1 _6793_ (.A1(_1807_),
    .A2(_1812_),
    .A3(_1850_),
    .B1(_1808_),
    .X(_1851_));
 sky130_fd_sc_hd__a21oi_1 _6794_ (.A1(_1800_),
    .A2(_1851_),
    .B1(_1801_),
    .Y(_1852_));
 sky130_fd_sc_hd__a221o_1 _6795_ (.A1(_1792_),
    .A2(_1795_),
    .B1(_1800_),
    .B2(_1851_),
    .C1(_1801_),
    .X(_1853_));
 sky130_fd_sc_hd__nand2_1 _6796_ (.A(_1796_),
    .B(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__a2bb2oi_1 _6797_ (.A1_N(_1788_),
    .A2_N(_1790_),
    .B1(_1796_),
    .B2(_1853_),
    .Y(_1855_));
 sky130_fd_sc_hd__and3_1 _6798_ (.A(_1708_),
    .B(_1709_),
    .C(_1710_),
    .X(_1856_));
 sky130_fd_sc_hd__a21oi_1 _6799_ (.A1(_1708_),
    .A2(_1709_),
    .B1(_1710_),
    .Y(_1857_));
 sky130_fd_sc_hd__or4_1 _6800_ (.A(_1791_),
    .B(_1855_),
    .C(_1856_),
    .D(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__o22a_1 _6801_ (.A1(_1791_),
    .A2(_1855_),
    .B1(_1856_),
    .B2(_1857_),
    .X(_1860_));
 sky130_fd_sc_hd__o22ai_1 _6802_ (.A1(_1791_),
    .A2(_1855_),
    .B1(_1856_),
    .B2(_1857_),
    .Y(_1861_));
 sky130_fd_sc_hd__and2_1 _6803_ (.A(net3),
    .B(net38),
    .X(_1862_));
 sky130_fd_sc_hd__o41a_1 _6804_ (.A1(_1791_),
    .A2(_1855_),
    .A3(_1856_),
    .A4(_1857_),
    .B1(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__or3_1 _6805_ (.A(_1786_),
    .B(_1860_),
    .C(_1863_),
    .X(_1864_));
 sky130_fd_sc_hd__a22o_2 _6806_ (.A1(_1778_),
    .A2(_1779_),
    .B1(_1785_),
    .B2(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__nand4_2 _6807_ (.A(_1778_),
    .B(_1779_),
    .C(_1785_),
    .D(_1864_),
    .Y(_1866_));
 sky130_fd_sc_hd__and2_1 _6808_ (.A(net5),
    .B(net38),
    .X(_1867_));
 sky130_fd_sc_hd__nand2_1 _6809_ (.A(net5),
    .B(net38),
    .Y(_1868_));
 sky130_fd_sc_hd__a41o_1 _6810_ (.A1(_1778_),
    .A2(_1779_),
    .A3(_1785_),
    .A4(_1864_),
    .B1(_1867_),
    .X(_1869_));
 sky130_fd_sc_hd__a31o_1 _6811_ (.A1(_1776_),
    .A2(_1865_),
    .A3(_1869_),
    .B1(_1777_),
    .X(_1871_));
 sky130_fd_sc_hd__xor2_1 _6812_ (.A(_1722_),
    .B(_1724_),
    .X(_1872_));
 sky130_fd_sc_hd__xnor2_1 _6813_ (.A(_1726_),
    .B(_1872_),
    .Y(_1873_));
 sky130_fd_sc_hd__and2_1 _6814_ (.A(_1871_),
    .B(_1873_),
    .X(_1874_));
 sky130_fd_sc_hd__nand2_1 _6815_ (.A(net7),
    .B(net38),
    .Y(_1875_));
 sky130_fd_sc_hd__o211a_1 _6816_ (.A1(_1871_),
    .A2(_1873_),
    .B1(net7),
    .C1(net38),
    .X(_1876_));
 sky130_fd_sc_hd__o31a_1 _6817_ (.A1(_1769_),
    .A2(_1874_),
    .A3(_1876_),
    .B1(_1768_),
    .X(_1877_));
 sky130_fd_sc_hd__xor2_1 _6818_ (.A(_1729_),
    .B(_1731_),
    .X(_1878_));
 sky130_fd_sc_hd__xnor2_2 _6819_ (.A(_1733_),
    .B(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hd__nor2_1 _6820_ (.A(_1877_),
    .B(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__nand2_1 _6821_ (.A(net9),
    .B(net38),
    .Y(_1882_));
 sky130_fd_sc_hd__a21boi_2 _6822_ (.A1(_1877_),
    .A2(_1879_),
    .B1_N(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__o31ai_4 _6823_ (.A1(_1762_),
    .A2(_1880_),
    .A3(_1883_),
    .B1(_1764_),
    .Y(_1884_));
 sky130_fd_sc_hd__xor2_1 _6824_ (.A(_1735_),
    .B(_1737_),
    .X(_1885_));
 sky130_fd_sc_hd__xnor2_1 _6825_ (.A(_1740_),
    .B(_1885_),
    .Y(_1886_));
 sky130_fd_sc_hd__or2_1 _6826_ (.A(_1884_),
    .B(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__nand2_1 _6827_ (.A(net11),
    .B(net38),
    .Y(_1888_));
 sky130_fd_sc_hd__a21bo_1 _6828_ (.A1(_1884_),
    .A2(_1886_),
    .B1_N(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__a31o_1 _6829_ (.A1(_1757_),
    .A2(_1887_),
    .A3(_1889_),
    .B1(_1755_),
    .X(_1890_));
 sky130_fd_sc_hd__xor2_1 _6830_ (.A(_1592_),
    .B(_1742_),
    .X(_1891_));
 sky130_fd_sc_hd__xnor2_2 _6831_ (.A(_1744_),
    .B(_1891_),
    .Y(_1893_));
 sky130_fd_sc_hd__nor2_1 _6832_ (.A(_1890_),
    .B(_1893_),
    .Y(_1894_));
 sky130_fd_sc_hd__nand2_1 _6833_ (.A(net14),
    .B(net38),
    .Y(_1895_));
 sky130_fd_sc_hd__a21boi_2 _6834_ (.A1(_1890_),
    .A2(_1893_),
    .B1_N(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__o31ai_2 _6835_ (.A1(_1748_),
    .A2(_1894_),
    .A3(_1896_),
    .B1(_1751_),
    .Y(_1897_));
 sky130_fd_sc_hd__a32o_1 _6836_ (.A1(_1589_),
    .A2(_1743_),
    .A3(_1745_),
    .B1(_1588_),
    .B2(net37),
    .X(_1898_));
 sky130_fd_sc_hd__and2_1 _6837_ (.A(net38),
    .B(_1716_),
    .X(_1899_));
 sky130_fd_sc_hd__o21ai_1 _6838_ (.A1(_1897_),
    .A2(_1898_),
    .B1(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__o21ai_1 _6839_ (.A1(_0088_),
    .A2(_1727_),
    .B1(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__nor2_1 _6840_ (.A(_0088_),
    .B(_1900_),
    .Y(_1902_));
 sky130_fd_sc_hd__o21ai_1 _6841_ (.A1(_0088_),
    .A2(_1900_),
    .B1(_1901_),
    .Y(_1904_));
 sky130_fd_sc_hd__xnor2_1 _6842_ (.A(_1897_),
    .B(_1898_),
    .Y(_1905_));
 sky130_fd_sc_hd__xnor2_1 _6843_ (.A(_1899_),
    .B(_1905_),
    .Y(_1906_));
 sky130_fd_sc_hd__o22ai_2 _6844_ (.A1(_1748_),
    .A2(_1750_),
    .B1(_1894_),
    .B2(_1896_),
    .Y(_1907_));
 sky130_fd_sc_hd__or4_1 _6845_ (.A(_1748_),
    .B(_1750_),
    .C(_1894_),
    .D(_1896_),
    .X(_1908_));
 sky130_fd_sc_hd__and4_1 _6846_ (.A(net14),
    .B(net39),
    .C(_1907_),
    .D(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__nand4_1 _6847_ (.A(net14),
    .B(net39),
    .C(_1907_),
    .D(_1908_),
    .Y(_1910_));
 sky130_fd_sc_hd__a22oi_2 _6848_ (.A1(net14),
    .A2(net39),
    .B1(_1907_),
    .B2(_1908_),
    .Y(_1911_));
 sky130_fd_sc_hd__xor2_1 _6849_ (.A(_1890_),
    .B(_1893_),
    .X(_1912_));
 sky130_fd_sc_hd__xnor2_1 _6850_ (.A(_1895_),
    .B(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__a22o_1 _6851_ (.A1(_1756_),
    .A2(_1757_),
    .B1(_1887_),
    .B2(_1889_),
    .X(_1915_));
 sky130_fd_sc_hd__nand4_2 _6852_ (.A(_1756_),
    .B(_1757_),
    .C(_1887_),
    .D(_1889_),
    .Y(_1916_));
 sky130_fd_sc_hd__and4_1 _6853_ (.A(net11),
    .B(net39),
    .C(_1915_),
    .D(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__a22oi_2 _6854_ (.A1(net11),
    .A2(net39),
    .B1(_1915_),
    .B2(_1916_),
    .Y(_1918_));
 sky130_fd_sc_hd__a22o_1 _6855_ (.A1(net11),
    .A2(net39),
    .B1(_1915_),
    .B2(_1916_),
    .X(_1919_));
 sky130_fd_sc_hd__o22ai_2 _6856_ (.A1(_1762_),
    .A2(_1763_),
    .B1(_1880_),
    .B2(_1883_),
    .Y(_1920_));
 sky130_fd_sc_hd__or4_1 _6857_ (.A(_1762_),
    .B(_1763_),
    .C(_1880_),
    .D(_1883_),
    .X(_1921_));
 sky130_fd_sc_hd__a22o_1 _6858_ (.A1(net9),
    .A2(net39),
    .B1(_1920_),
    .B2(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__and4_1 _6859_ (.A(net9),
    .B(net39),
    .C(_1920_),
    .D(_1921_),
    .X(_1923_));
 sky130_fd_sc_hd__nand4_1 _6860_ (.A(net9),
    .B(net39),
    .C(_1920_),
    .D(_1921_),
    .Y(_1924_));
 sky130_fd_sc_hd__and2_1 _6861_ (.A(net7),
    .B(net39),
    .X(_1926_));
 sky130_fd_sc_hd__o211ai_2 _6862_ (.A1(_1874_),
    .A2(_1876_),
    .B1(_1768_),
    .C1(_1770_),
    .Y(_1927_));
 sky130_fd_sc_hd__a211o_1 _6863_ (.A1(_1768_),
    .A2(_1770_),
    .B1(_1874_),
    .C1(_1876_),
    .X(_1928_));
 sky130_fd_sc_hd__a21oi_1 _6864_ (.A1(_1927_),
    .A2(_1928_),
    .B1(_1926_),
    .Y(_1929_));
 sky130_fd_sc_hd__a21o_1 _6865_ (.A1(_1927_),
    .A2(_1928_),
    .B1(_1926_),
    .X(_1930_));
 sky130_fd_sc_hd__and3_1 _6866_ (.A(_1926_),
    .B(_1927_),
    .C(_1928_),
    .X(_1931_));
 sky130_fd_sc_hd__nand2_1 _6867_ (.A(net5),
    .B(net39),
    .Y(_1932_));
 sky130_fd_sc_hd__o211ai_2 _6868_ (.A1(_1775_),
    .A2(_1777_),
    .B1(_1865_),
    .C1(_1869_),
    .Y(_1933_));
 sky130_fd_sc_hd__a211o_1 _6869_ (.A1(_1865_),
    .A2(_1869_),
    .B1(_1775_),
    .C1(_1777_),
    .X(_1934_));
 sky130_fd_sc_hd__a21oi_1 _6870_ (.A1(_1933_),
    .A2(_1934_),
    .B1(_1932_),
    .Y(_1935_));
 sky130_fd_sc_hd__a21o_1 _6871_ (.A1(_1933_),
    .A2(_1934_),
    .B1(_1932_),
    .X(_1937_));
 sky130_fd_sc_hd__and3_1 _6872_ (.A(_1932_),
    .B(_1933_),
    .C(_1934_),
    .X(_1938_));
 sky130_fd_sc_hd__nand2_1 _6873_ (.A(net3),
    .B(net39),
    .Y(_1939_));
 sky130_fd_sc_hd__o22ai_1 _6874_ (.A1(_1784_),
    .A2(_1786_),
    .B1(_1860_),
    .B2(_1863_),
    .Y(_1940_));
 sky130_fd_sc_hd__or4_1 _6875_ (.A(_1784_),
    .B(_1786_),
    .C(_1860_),
    .D(_1863_),
    .X(_1941_));
 sky130_fd_sc_hd__a21o_1 _6876_ (.A1(_1940_),
    .A2(_1941_),
    .B1(_1939_),
    .X(_1942_));
 sky130_fd_sc_hd__nand3_1 _6877_ (.A(_1939_),
    .B(_1940_),
    .C(_1941_),
    .Y(_1943_));
 sky130_fd_sc_hd__nand2_1 _6878_ (.A(net32),
    .B(net39),
    .Y(_1944_));
 sky130_fd_sc_hd__inv_2 _6879_ (.A(_1944_),
    .Y(_1945_));
 sky130_fd_sc_hd__xnor2_1 _6880_ (.A(_1788_),
    .B(_1790_),
    .Y(_1946_));
 sky130_fd_sc_hd__xnor2_1 _6881_ (.A(_1854_),
    .B(_1946_),
    .Y(_1948_));
 sky130_fd_sc_hd__or2_1 _6882_ (.A(_1945_),
    .B(_1948_),
    .X(_1949_));
 sky130_fd_sc_hd__nand2_1 _6883_ (.A(net31),
    .B(net39),
    .Y(_1950_));
 sky130_fd_sc_hd__xnor2_1 _6884_ (.A(_1792_),
    .B(_1795_),
    .Y(_1951_));
 sky130_fd_sc_hd__xnor2_1 _6885_ (.A(_1852_),
    .B(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__nand2b_1 _6886_ (.A_N(_1952_),
    .B(_1950_),
    .Y(_1953_));
 sky130_fd_sc_hd__and3_1 _6887_ (.A(net31),
    .B(net39),
    .C(_1952_),
    .X(_1954_));
 sky130_fd_sc_hd__nand2_1 _6888_ (.A(net30),
    .B(net39),
    .Y(_1955_));
 sky130_fd_sc_hd__xnor2_1 _6889_ (.A(_1797_),
    .B(_1799_),
    .Y(_1956_));
 sky130_fd_sc_hd__xnor2_1 _6890_ (.A(_1851_),
    .B(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__a21o_1 _6891_ (.A1(net30),
    .A2(net39),
    .B1(_1957_),
    .X(_1959_));
 sky130_fd_sc_hd__and3_1 _6892_ (.A(net30),
    .B(net39),
    .C(_1957_),
    .X(_1960_));
 sky130_fd_sc_hd__and2_1 _6893_ (.A(net29),
    .B(net39),
    .X(_1961_));
 sky130_fd_sc_hd__o211ai_2 _6894_ (.A1(_1806_),
    .A2(_1808_),
    .B1(_1812_),
    .C1(_1850_),
    .Y(_1962_));
 sky130_fd_sc_hd__a211o_1 _6895_ (.A1(_1812_),
    .A2(_1850_),
    .B1(_1806_),
    .C1(_1808_),
    .X(_1963_));
 sky130_fd_sc_hd__and3_1 _6896_ (.A(_1961_),
    .B(_1962_),
    .C(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__a21oi_1 _6897_ (.A1(_1962_),
    .A2(_1963_),
    .B1(_1961_),
    .Y(_1965_));
 sky130_fd_sc_hd__a21o_1 _6898_ (.A1(_1962_),
    .A2(_1963_),
    .B1(_1961_),
    .X(_1966_));
 sky130_fd_sc_hd__nand2_1 _6899_ (.A(net28),
    .B(net39),
    .Y(_1967_));
 sky130_fd_sc_hd__inv_2 _6900_ (.A(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__xnor2_1 _6901_ (.A(_1809_),
    .B(_1811_),
    .Y(_1970_));
 sky130_fd_sc_hd__xnor2_1 _6902_ (.A(_1849_),
    .B(_1970_),
    .Y(_1971_));
 sky130_fd_sc_hd__or2_1 _6903_ (.A(_1968_),
    .B(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__xnor2_1 _6904_ (.A(_1813_),
    .B(_1817_),
    .Y(_1973_));
 sky130_fd_sc_hd__xnor2_1 _6905_ (.A(_1846_),
    .B(_1973_),
    .Y(_1974_));
 sky130_fd_sc_hd__nand2_1 _6906_ (.A(net27),
    .B(net39),
    .Y(_1975_));
 sky130_fd_sc_hd__and3_1 _6907_ (.A(net27),
    .B(net39),
    .C(_1974_),
    .X(_1976_));
 sky130_fd_sc_hd__nand2b_1 _6908_ (.A_N(_1974_),
    .B(_1975_),
    .Y(_1977_));
 sky130_fd_sc_hd__nand2_1 _6909_ (.A(net26),
    .B(net39),
    .Y(_1978_));
 sky130_fd_sc_hd__xor2_1 _6910_ (.A(_1819_),
    .B(_1821_),
    .X(_1979_));
 sky130_fd_sc_hd__xnor2_1 _6911_ (.A(_1845_),
    .B(_1979_),
    .Y(_1981_));
 sky130_fd_sc_hd__a21o_1 _6912_ (.A1(net26),
    .A2(net39),
    .B1(_1981_),
    .X(_1982_));
 sky130_fd_sc_hd__and3_1 _6913_ (.A(net26),
    .B(net39),
    .C(_1981_),
    .X(_1983_));
 sky130_fd_sc_hd__a21o_1 _6914_ (.A1(_1827_),
    .A2(_1828_),
    .B1(_1844_),
    .X(_1984_));
 sky130_fd_sc_hd__nand3_1 _6915_ (.A(_1827_),
    .B(_1828_),
    .C(_1844_),
    .Y(_1985_));
 sky130_fd_sc_hd__a22o_1 _6916_ (.A1(net23),
    .A2(net39),
    .B1(_1984_),
    .B2(_1985_),
    .X(_1986_));
 sky130_fd_sc_hd__nand4_1 _6917_ (.A(net23),
    .B(net39),
    .C(_1984_),
    .D(_1985_),
    .Y(_1987_));
 sky130_fd_sc_hd__or4bb_1 _6918_ (.A(_1832_),
    .B(_1834_),
    .C_N(_1839_),
    .D_N(_1843_),
    .X(_1988_));
 sky130_fd_sc_hd__a2bb2o_1 _6919_ (.A1_N(_1832_),
    .A2_N(_1834_),
    .B1(_1839_),
    .B2(_1843_),
    .X(_1989_));
 sky130_fd_sc_hd__nand2_1 _6920_ (.A(net12),
    .B(net39),
    .Y(_1990_));
 sky130_fd_sc_hd__and3_1 _6921_ (.A(_1988_),
    .B(_1989_),
    .C(_1990_),
    .X(_1992_));
 sky130_fd_sc_hd__a21o_1 _6922_ (.A1(_1988_),
    .A2(_1989_),
    .B1(_1990_),
    .X(_1993_));
 sky130_fd_sc_hd__xnor2_1 _6923_ (.A(_1835_),
    .B(_1838_),
    .Y(_1994_));
 sky130_fd_sc_hd__xor2_1 _6924_ (.A(_1842_),
    .B(_1994_),
    .X(_1995_));
 sky130_fd_sc_hd__or3b_1 _6925_ (.A(_4198_),
    .B(_0088_),
    .C_N(_1995_),
    .X(_1996_));
 sky130_fd_sc_hd__o21ai_1 _6926_ (.A1(_1992_),
    .A2(_1996_),
    .B1(_1993_),
    .Y(_1997_));
 sky130_fd_sc_hd__o21a_1 _6927_ (.A1(_1992_),
    .A2(_1996_),
    .B1(_1993_),
    .X(_1998_));
 sky130_fd_sc_hd__a21bo_1 _6928_ (.A1(_1986_),
    .A2(_1997_),
    .B1_N(_1987_),
    .X(_1999_));
 sky130_fd_sc_hd__a21o_1 _6929_ (.A1(_1982_),
    .A2(_1999_),
    .B1(_1983_),
    .X(_2000_));
 sky130_fd_sc_hd__a21oi_1 _6930_ (.A1(_1977_),
    .A2(_2000_),
    .B1(_1976_),
    .Y(_2001_));
 sky130_fd_sc_hd__a221o_1 _6931_ (.A1(_1968_),
    .A2(_1971_),
    .B1(_1977_),
    .B2(_2000_),
    .C1(_1976_),
    .X(_2003_));
 sky130_fd_sc_hd__a21o_1 _6932_ (.A1(_1972_),
    .A2(_2003_),
    .B1(_1964_),
    .X(_2004_));
 sky130_fd_sc_hd__a31o_1 _6933_ (.A1(_1959_),
    .A2(_1966_),
    .A3(_2004_),
    .B1(_1960_),
    .X(_2005_));
 sky130_fd_sc_hd__a21oi_1 _6934_ (.A1(_1953_),
    .A2(_2005_),
    .B1(_1954_),
    .Y(_2006_));
 sky130_fd_sc_hd__a221o_1 _6935_ (.A1(_1945_),
    .A2(_1948_),
    .B1(_1953_),
    .B2(_2005_),
    .C1(_1954_),
    .X(_2007_));
 sky130_fd_sc_hd__a21o_1 _6936_ (.A1(_1858_),
    .A2(_1861_),
    .B1(_1862_),
    .X(_2008_));
 sky130_fd_sc_hd__nand3_1 _6937_ (.A(_1858_),
    .B(_1861_),
    .C(_1862_),
    .Y(_2009_));
 sky130_fd_sc_hd__a22o_1 _6938_ (.A1(_1949_),
    .A2(_2007_),
    .B1(_2008_),
    .B2(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__nand4_2 _6939_ (.A(_1949_),
    .B(_2007_),
    .C(_2008_),
    .D(_2009_),
    .Y(_2011_));
 sky130_fd_sc_hd__and2_1 _6940_ (.A(net2),
    .B(net39),
    .X(_2012_));
 sky130_fd_sc_hd__nand2_1 _6941_ (.A(net2),
    .B(net39),
    .Y(_2014_));
 sky130_fd_sc_hd__a41o_1 _6942_ (.A1(_1949_),
    .A2(_2007_),
    .A3(_2008_),
    .A4(_2009_),
    .B1(_2012_),
    .X(_2015_));
 sky130_fd_sc_hd__nand3_1 _6943_ (.A(_1943_),
    .B(_2010_),
    .C(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__nand3_1 _6944_ (.A(_1865_),
    .B(_1866_),
    .C(_1868_),
    .Y(_2017_));
 sky130_fd_sc_hd__a21o_1 _6945_ (.A1(_1865_),
    .A2(_1866_),
    .B1(_1868_),
    .X(_2018_));
 sky130_fd_sc_hd__a21oi_1 _6946_ (.A1(_1865_),
    .A2(_1866_),
    .B1(_1867_),
    .Y(_2019_));
 sky130_fd_sc_hd__and3_1 _6947_ (.A(_1865_),
    .B(_1866_),
    .C(_1867_),
    .X(_2020_));
 sky130_fd_sc_hd__o211ai_1 _6948_ (.A1(_2019_),
    .A2(_2020_),
    .B1(_1942_),
    .C1(_2016_),
    .Y(_2021_));
 sky130_fd_sc_hd__a211o_1 _6949_ (.A1(_1942_),
    .A2(_2016_),
    .B1(_2019_),
    .C1(_2020_),
    .X(_2022_));
 sky130_fd_sc_hd__nand2_1 _6950_ (.A(net4),
    .B(net39),
    .Y(_2023_));
 sky130_fd_sc_hd__a41o_1 _6951_ (.A1(_1942_),
    .A2(_2016_),
    .A3(_2017_),
    .A4(_2018_),
    .B1(_2023_),
    .X(_2025_));
 sky130_fd_sc_hd__a31o_1 _6952_ (.A1(_1937_),
    .A2(_2022_),
    .A3(_2025_),
    .B1(_1938_),
    .X(_2026_));
 sky130_fd_sc_hd__xnor2_1 _6953_ (.A(_1871_),
    .B(_1873_),
    .Y(_2027_));
 sky130_fd_sc_hd__xnor2_2 _6954_ (.A(_1875_),
    .B(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__nand2_1 _6955_ (.A(_2026_),
    .B(_2028_),
    .Y(_2029_));
 sky130_fd_sc_hd__and2_1 _6956_ (.A(net6),
    .B(net39),
    .X(_2030_));
 sky130_fd_sc_hd__o21bai_2 _6957_ (.A1(_2026_),
    .A2(_2028_),
    .B1_N(_2030_),
    .Y(_2031_));
 sky130_fd_sc_hd__a31o_1 _6958_ (.A1(_1930_),
    .A2(_2029_),
    .A3(_2031_),
    .B1(_1931_),
    .X(_2032_));
 sky130_fd_sc_hd__xor2_1 _6959_ (.A(_1877_),
    .B(_1879_),
    .X(_2033_));
 sky130_fd_sc_hd__xnor2_1 _6960_ (.A(_1882_),
    .B(_2033_),
    .Y(_2034_));
 sky130_fd_sc_hd__or2_1 _6961_ (.A(_2032_),
    .B(_2034_),
    .X(_2036_));
 sky130_fd_sc_hd__nand2_1 _6962_ (.A(net8),
    .B(net39),
    .Y(_2037_));
 sky130_fd_sc_hd__a21bo_1 _6963_ (.A1(_2032_),
    .A2(_2034_),
    .B1_N(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__a31o_1 _6964_ (.A1(_1922_),
    .A2(_2036_),
    .A3(_2038_),
    .B1(_1923_),
    .X(_2039_));
 sky130_fd_sc_hd__xor2_1 _6965_ (.A(_1884_),
    .B(_1886_),
    .X(_2040_));
 sky130_fd_sc_hd__xnor2_1 _6966_ (.A(_1888_),
    .B(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__or2_1 _6967_ (.A(_2039_),
    .B(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__nand2_1 _6968_ (.A(net10),
    .B(net39),
    .Y(_2043_));
 sky130_fd_sc_hd__a21bo_1 _6969_ (.A1(_2039_),
    .A2(_2041_),
    .B1_N(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__a31o_1 _6970_ (.A1(_1919_),
    .A2(_2042_),
    .A3(_2044_),
    .B1(_1917_),
    .X(_2045_));
 sky130_fd_sc_hd__nor2_1 _6971_ (.A(_1913_),
    .B(_2045_),
    .Y(_2047_));
 sky130_fd_sc_hd__nor2_1 _6972_ (.A(_0000_),
    .B(_0088_),
    .Y(_2048_));
 sky130_fd_sc_hd__a21oi_1 _6973_ (.A1(_1913_),
    .A2(_2045_),
    .B1(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__o31ai_2 _6974_ (.A1(_1911_),
    .A2(_2047_),
    .A3(_2049_),
    .B1(_1910_),
    .Y(_2050_));
 sky130_fd_sc_hd__or2_1 _6975_ (.A(_1906_),
    .B(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__nand2_1 _6976_ (.A(net15),
    .B(net39),
    .Y(_2052_));
 sky130_fd_sc_hd__a21bo_1 _6977_ (.A1(_1906_),
    .A2(_2050_),
    .B1_N(_2052_),
    .X(_2053_));
 sky130_fd_sc_hd__nand3_1 _6978_ (.A(_1904_),
    .B(_2051_),
    .C(_2053_),
    .Y(_2054_));
 sky130_fd_sc_hd__a21o_1 _6979_ (.A1(_2051_),
    .A2(_2053_),
    .B1(_1904_),
    .X(_2055_));
 sky130_fd_sc_hd__a21oi_2 _6980_ (.A1(_2054_),
    .A2(_2055_),
    .B1(_3979_),
    .Y(_2056_));
 sky130_fd_sc_hd__and3_1 _6981_ (.A(_3979_),
    .B(_2054_),
    .C(_2055_),
    .X(_2058_));
 sky130_fd_sc_hd__nand3_1 _6982_ (.A(_3979_),
    .B(_2054_),
    .C(_2055_),
    .Y(_2059_));
 sky130_fd_sc_hd__nor2_1 _6983_ (.A(_0000_),
    .B(_0099_),
    .Y(_2060_));
 sky130_fd_sc_hd__o22ai_1 _6984_ (.A1(_1909_),
    .A2(_1911_),
    .B1(_2047_),
    .B2(_2049_),
    .Y(_2061_));
 sky130_fd_sc_hd__or4_1 _6985_ (.A(_1909_),
    .B(_1911_),
    .C(_2047_),
    .D(_2049_),
    .X(_2062_));
 sky130_fd_sc_hd__a21oi_1 _6986_ (.A1(_2061_),
    .A2(_2062_),
    .B1(_2060_),
    .Y(_2063_));
 sky130_fd_sc_hd__and3_1 _6987_ (.A(_2060_),
    .B(_2061_),
    .C(_2062_),
    .X(_2064_));
 sky130_fd_sc_hd__nand3_1 _6988_ (.A(_2060_),
    .B(_2061_),
    .C(_2062_),
    .Y(_2065_));
 sky130_fd_sc_hd__nand2_1 _6989_ (.A(net10),
    .B(net40),
    .Y(_2066_));
 sky130_fd_sc_hd__o211ai_2 _6990_ (.A1(_1917_),
    .A2(_1918_),
    .B1(_2042_),
    .C1(_2044_),
    .Y(_2067_));
 sky130_fd_sc_hd__a211o_1 _6991_ (.A1(_2042_),
    .A2(_2044_),
    .B1(_1917_),
    .C1(_1918_),
    .X(_2069_));
 sky130_fd_sc_hd__and3_1 _6992_ (.A(_2066_),
    .B(_2067_),
    .C(_2069_),
    .X(_2070_));
 sky130_fd_sc_hd__nand3_1 _6993_ (.A(_2066_),
    .B(_2067_),
    .C(_2069_),
    .Y(_2071_));
 sky130_fd_sc_hd__a21oi_1 _6994_ (.A1(_2067_),
    .A2(_2069_),
    .B1(_2066_),
    .Y(_2072_));
 sky130_fd_sc_hd__and2_1 _6995_ (.A(net8),
    .B(net40),
    .X(_2073_));
 sky130_fd_sc_hd__a22o_1 _6996_ (.A1(_1922_),
    .A2(_1924_),
    .B1(_2036_),
    .B2(_2038_),
    .X(_2074_));
 sky130_fd_sc_hd__nand4_1 _6997_ (.A(_1922_),
    .B(_1924_),
    .C(_2036_),
    .D(_2038_),
    .Y(_2075_));
 sky130_fd_sc_hd__a21oi_1 _6998_ (.A1(_2074_),
    .A2(_2075_),
    .B1(_2073_),
    .Y(_2076_));
 sky130_fd_sc_hd__a21o_1 _6999_ (.A1(_2074_),
    .A2(_2075_),
    .B1(_2073_),
    .X(_2077_));
 sky130_fd_sc_hd__and3_1 _7000_ (.A(_2073_),
    .B(_2074_),
    .C(_2075_),
    .X(_2078_));
 sky130_fd_sc_hd__nand2_1 _7001_ (.A(net6),
    .B(net40),
    .Y(_2080_));
 sky130_fd_sc_hd__o211ai_2 _7002_ (.A1(_1929_),
    .A2(_1931_),
    .B1(_2029_),
    .C1(_2031_),
    .Y(_2081_));
 sky130_fd_sc_hd__a211o_1 _7003_ (.A1(_2029_),
    .A2(_2031_),
    .B1(_1929_),
    .C1(_1931_),
    .X(_2082_));
 sky130_fd_sc_hd__a21oi_1 _7004_ (.A1(_2081_),
    .A2(_2082_),
    .B1(_2080_),
    .Y(_2083_));
 sky130_fd_sc_hd__a21o_1 _7005_ (.A1(_2081_),
    .A2(_2082_),
    .B1(_2080_),
    .X(_2084_));
 sky130_fd_sc_hd__and3_1 _7006_ (.A(_2080_),
    .B(_2081_),
    .C(_2082_),
    .X(_2085_));
 sky130_fd_sc_hd__and2_1 _7007_ (.A(net4),
    .B(net40),
    .X(_2086_));
 sky130_fd_sc_hd__o211ai_2 _7008_ (.A1(_1935_),
    .A2(_1938_),
    .B1(_2022_),
    .C1(_2025_),
    .Y(_2087_));
 sky130_fd_sc_hd__a211o_1 _7009_ (.A1(_2022_),
    .A2(_2025_),
    .B1(_1935_),
    .C1(_1938_),
    .X(_2088_));
 sky130_fd_sc_hd__a21oi_1 _7010_ (.A1(_2087_),
    .A2(_2088_),
    .B1(_2086_),
    .Y(_2089_));
 sky130_fd_sc_hd__and3_1 _7011_ (.A(_2086_),
    .B(_2087_),
    .C(_2088_),
    .X(_2091_));
 sky130_fd_sc_hd__nand3_1 _7012_ (.A(_2086_),
    .B(_2087_),
    .C(_2088_),
    .Y(_2092_));
 sky130_fd_sc_hd__and2_1 _7013_ (.A(net2),
    .B(net40),
    .X(_2093_));
 sky130_fd_sc_hd__a22o_1 _7014_ (.A1(_1942_),
    .A2(_1943_),
    .B1(_2010_),
    .B2(_2015_),
    .X(_2094_));
 sky130_fd_sc_hd__nand4_1 _7015_ (.A(_1942_),
    .B(_1943_),
    .C(_2010_),
    .D(_2015_),
    .Y(_2095_));
 sky130_fd_sc_hd__a21o_1 _7016_ (.A1(_2094_),
    .A2(_2095_),
    .B1(_2093_),
    .X(_2096_));
 sky130_fd_sc_hd__and3_1 _7017_ (.A(_2093_),
    .B(_2094_),
    .C(_2095_),
    .X(_2097_));
 sky130_fd_sc_hd__nand3_1 _7018_ (.A(_2093_),
    .B(_2094_),
    .C(_2095_),
    .Y(_2098_));
 sky130_fd_sc_hd__xnor2_1 _7019_ (.A(_1944_),
    .B(_1948_),
    .Y(_2099_));
 sky130_fd_sc_hd__xnor2_1 _7020_ (.A(_2006_),
    .B(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__and2_1 _7021_ (.A(net31),
    .B(net40),
    .X(_2102_));
 sky130_fd_sc_hd__or2_1 _7022_ (.A(_2100_),
    .B(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__and2_1 _7023_ (.A(net30),
    .B(net40),
    .X(_2104_));
 sky130_fd_sc_hd__xor2_1 _7024_ (.A(_1950_),
    .B(_1952_),
    .X(_2105_));
 sky130_fd_sc_hd__xnor2_1 _7025_ (.A(_2005_),
    .B(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__and2_1 _7026_ (.A(_2104_),
    .B(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__xnor2_1 _7027_ (.A(_1955_),
    .B(_1957_),
    .Y(_2108_));
 sky130_fd_sc_hd__a21o_1 _7028_ (.A1(_1966_),
    .A2(_2004_),
    .B1(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__nand3_1 _7029_ (.A(_1966_),
    .B(_2004_),
    .C(_2108_),
    .Y(_2110_));
 sky130_fd_sc_hd__and4_1 _7030_ (.A(net29),
    .B(net40),
    .C(_2109_),
    .D(_2110_),
    .X(_2111_));
 sky130_fd_sc_hd__a22oi_1 _7031_ (.A1(net29),
    .A2(net40),
    .B1(_2109_),
    .B2(_2110_),
    .Y(_2113_));
 sky130_fd_sc_hd__a22o_1 _7032_ (.A1(net29),
    .A2(net40),
    .B1(_2109_),
    .B2(_2110_),
    .X(_2114_));
 sky130_fd_sc_hd__and2_1 _7033_ (.A(net28),
    .B(net40),
    .X(_2115_));
 sky130_fd_sc_hd__a2bb2o_1 _7034_ (.A1_N(_1964_),
    .A2_N(_1965_),
    .B1(_1972_),
    .B2(_2003_),
    .X(_2116_));
 sky130_fd_sc_hd__or4bb_1 _7035_ (.A(_1964_),
    .B(_1965_),
    .C_N(_1972_),
    .D_N(_2003_),
    .X(_2117_));
 sky130_fd_sc_hd__a21o_1 _7036_ (.A1(_2116_),
    .A2(_2117_),
    .B1(_2115_),
    .X(_2118_));
 sky130_fd_sc_hd__and3_1 _7037_ (.A(_2115_),
    .B(_2116_),
    .C(_2117_),
    .X(_2119_));
 sky130_fd_sc_hd__nand3_1 _7038_ (.A(_2115_),
    .B(_2116_),
    .C(_2117_),
    .Y(_2120_));
 sky130_fd_sc_hd__nor2_1 _7039_ (.A(_4187_),
    .B(_0099_),
    .Y(_2121_));
 sky130_fd_sc_hd__xnor2_1 _7040_ (.A(_1967_),
    .B(_1971_),
    .Y(_2122_));
 sky130_fd_sc_hd__xnor2_1 _7041_ (.A(_2001_),
    .B(_2122_),
    .Y(_2124_));
 sky130_fd_sc_hd__or2_1 _7042_ (.A(_2121_),
    .B(_2124_),
    .X(_2125_));
 sky130_fd_sc_hd__nand2_1 _7043_ (.A(net26),
    .B(net40),
    .Y(_2126_));
 sky130_fd_sc_hd__xor2_1 _7044_ (.A(_1974_),
    .B(_1975_),
    .X(_2127_));
 sky130_fd_sc_hd__xnor2_1 _7045_ (.A(_2000_),
    .B(_2127_),
    .Y(_2128_));
 sky130_fd_sc_hd__a21o_1 _7046_ (.A1(net26),
    .A2(net40),
    .B1(_2128_),
    .X(_2129_));
 sky130_fd_sc_hd__and2_1 _7047_ (.A(net23),
    .B(net40),
    .X(_2130_));
 sky130_fd_sc_hd__xor2_1 _7048_ (.A(_1978_),
    .B(_1981_),
    .X(_2131_));
 sky130_fd_sc_hd__xnor2_1 _7049_ (.A(_1999_),
    .B(_2131_),
    .Y(_2132_));
 sky130_fd_sc_hd__and2_1 _7050_ (.A(_2130_),
    .B(_2132_),
    .X(_2133_));
 sky130_fd_sc_hd__nand2_1 _7051_ (.A(net12),
    .B(net40),
    .Y(_2135_));
 sky130_fd_sc_hd__a21o_1 _7052_ (.A1(_1986_),
    .A2(_1987_),
    .B1(_1998_),
    .X(_2136_));
 sky130_fd_sc_hd__nand3_1 _7053_ (.A(_1986_),
    .B(_1987_),
    .C(_1998_),
    .Y(_2137_));
 sky130_fd_sc_hd__a21o_1 _7054_ (.A1(_2136_),
    .A2(_2137_),
    .B1(_2135_),
    .X(_2138_));
 sky130_fd_sc_hd__or2_1 _7055_ (.A(_1993_),
    .B(_1996_),
    .X(_2139_));
 sky130_fd_sc_hd__nand2_1 _7056_ (.A(net1),
    .B(net40),
    .Y(_2140_));
 sky130_fd_sc_hd__a221o_1 _7057_ (.A1(_1992_),
    .A2(_1996_),
    .B1(_1997_),
    .B2(_2139_),
    .C1(_2140_),
    .X(_2141_));
 sky130_fd_sc_hd__a31o_1 _7058_ (.A1(_2135_),
    .A2(_2136_),
    .A3(_2137_),
    .B1(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__nand2_1 _7059_ (.A(_2138_),
    .B(_2142_),
    .Y(_2143_));
 sky130_fd_sc_hd__o2bb2a_1 _7060_ (.A1_N(_2138_),
    .A2_N(_2142_),
    .B1(_2130_),
    .B2(_2132_),
    .X(_2144_));
 sky130_fd_sc_hd__or2_1 _7061_ (.A(_2133_),
    .B(_2144_),
    .X(_2146_));
 sky130_fd_sc_hd__a311o_1 _7062_ (.A1(net26),
    .A2(net40),
    .A3(_2128_),
    .B1(_2133_),
    .C1(_2144_),
    .X(_2147_));
 sky130_fd_sc_hd__and2_1 _7063_ (.A(_2129_),
    .B(_2147_),
    .X(_2148_));
 sky130_fd_sc_hd__a22o_1 _7064_ (.A1(_2121_),
    .A2(_2124_),
    .B1(_2129_),
    .B2(_2147_),
    .X(_2149_));
 sky130_fd_sc_hd__a31o_1 _7065_ (.A1(_2118_),
    .A2(_2125_),
    .A3(_2149_),
    .B1(_2119_),
    .X(_2150_));
 sky130_fd_sc_hd__o21a_1 _7066_ (.A1(_2111_),
    .A2(_2150_),
    .B1(_2114_),
    .X(_2151_));
 sky130_fd_sc_hd__o221a_1 _7067_ (.A1(_2104_),
    .A2(_2106_),
    .B1(_2111_),
    .B2(_2150_),
    .C1(_2114_),
    .X(_2152_));
 sky130_fd_sc_hd__or2_1 _7068_ (.A(_2107_),
    .B(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__a211o_1 _7069_ (.A1(_2100_),
    .A2(_2102_),
    .B1(_2107_),
    .C1(_2152_),
    .X(_2154_));
 sky130_fd_sc_hd__and3_1 _7070_ (.A(_2010_),
    .B(_2011_),
    .C(_2014_),
    .X(_2155_));
 sky130_fd_sc_hd__a21oi_1 _7071_ (.A1(_2010_),
    .A2(_2011_),
    .B1(_2014_),
    .Y(_2157_));
 sky130_fd_sc_hd__a21o_1 _7072_ (.A1(_2010_),
    .A2(_2011_),
    .B1(_2012_),
    .X(_2158_));
 sky130_fd_sc_hd__nand4_1 _7073_ (.A(net2),
    .B(net39),
    .C(_2010_),
    .D(_2011_),
    .Y(_2159_));
 sky130_fd_sc_hd__a211o_1 _7074_ (.A1(_2103_),
    .A2(_2154_),
    .B1(_2155_),
    .C1(_2157_),
    .X(_2160_));
 sky130_fd_sc_hd__o211ai_1 _7075_ (.A1(_2155_),
    .A2(_2157_),
    .B1(_2103_),
    .C1(_2154_),
    .Y(_2161_));
 sky130_fd_sc_hd__and2_1 _7076_ (.A(net32),
    .B(net40),
    .X(_2162_));
 sky130_fd_sc_hd__a41o_1 _7077_ (.A1(_2103_),
    .A2(_2154_),
    .A3(_2158_),
    .A4(_2159_),
    .B1(_2162_),
    .X(_2163_));
 sky130_fd_sc_hd__a31oi_2 _7078_ (.A1(_2096_),
    .A2(_2160_),
    .A3(_2163_),
    .B1(_2097_),
    .Y(_2164_));
 sky130_fd_sc_hd__nand3_1 _7079_ (.A(_2021_),
    .B(_2022_),
    .C(_2023_),
    .Y(_2165_));
 sky130_fd_sc_hd__a21o_1 _7080_ (.A1(_2021_),
    .A2(_2022_),
    .B1(_2023_),
    .X(_2166_));
 sky130_fd_sc_hd__nand3_1 _7081_ (.A(_2164_),
    .B(_2165_),
    .C(_2166_),
    .Y(_2168_));
 sky130_fd_sc_hd__a21o_1 _7082_ (.A1(_2165_),
    .A2(_2166_),
    .B1(_2164_),
    .X(_2169_));
 sky130_fd_sc_hd__nor2_1 _7083_ (.A(_0011_),
    .B(_0099_),
    .Y(_2170_));
 sky130_fd_sc_hd__a311o_1 _7084_ (.A1(_2164_),
    .A2(_2165_),
    .A3(_2166_),
    .B1(_0099_),
    .C1(_0011_),
    .X(_2171_));
 sky130_fd_sc_hd__a31oi_2 _7085_ (.A1(_2092_),
    .A2(_2169_),
    .A3(_2171_),
    .B1(_2089_),
    .Y(_2172_));
 sky130_fd_sc_hd__xnor2_1 _7086_ (.A(_2026_),
    .B(_2028_),
    .Y(_2173_));
 sky130_fd_sc_hd__xnor2_2 _7087_ (.A(_2030_),
    .B(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__nand2_1 _7088_ (.A(_2172_),
    .B(_2174_),
    .Y(_2175_));
 sky130_fd_sc_hd__nand2_1 _7089_ (.A(net5),
    .B(net40),
    .Y(_2176_));
 sky130_fd_sc_hd__o211ai_2 _7090_ (.A1(_2172_),
    .A2(_2174_),
    .B1(net5),
    .C1(net40),
    .Y(_2177_));
 sky130_fd_sc_hd__a31oi_2 _7091_ (.A1(_2084_),
    .A2(_2175_),
    .A3(_2177_),
    .B1(_2085_),
    .Y(_2179_));
 sky130_fd_sc_hd__xor2_1 _7092_ (.A(_2032_),
    .B(_2034_),
    .X(_2180_));
 sky130_fd_sc_hd__xnor2_1 _7093_ (.A(_2037_),
    .B(_2180_),
    .Y(_2181_));
 sky130_fd_sc_hd__or2_1 _7094_ (.A(_2179_),
    .B(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__nand2_1 _7095_ (.A(net7),
    .B(net40),
    .Y(_2183_));
 sky130_fd_sc_hd__a21bo_1 _7096_ (.A1(_2179_),
    .A2(_2181_),
    .B1_N(_2183_),
    .X(_2184_));
 sky130_fd_sc_hd__a31o_1 _7097_ (.A1(_2077_),
    .A2(_2182_),
    .A3(_2184_),
    .B1(_2078_),
    .X(_2185_));
 sky130_fd_sc_hd__xor2_1 _7098_ (.A(_2039_),
    .B(_2041_),
    .X(_2186_));
 sky130_fd_sc_hd__xnor2_1 _7099_ (.A(_2043_),
    .B(_2186_),
    .Y(_2187_));
 sky130_fd_sc_hd__or2_1 _7100_ (.A(_2185_),
    .B(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__nand2_1 _7101_ (.A(net9),
    .B(net40),
    .Y(_2190_));
 sky130_fd_sc_hd__a21bo_1 _7102_ (.A1(_2185_),
    .A2(_2187_),
    .B1_N(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__a31o_1 _7103_ (.A1(_2071_),
    .A2(_2188_),
    .A3(_2191_),
    .B1(_2072_),
    .X(_2192_));
 sky130_fd_sc_hd__xnor2_1 _7104_ (.A(_1913_),
    .B(_2045_),
    .Y(_2193_));
 sky130_fd_sc_hd__xnor2_1 _7105_ (.A(_2048_),
    .B(_2193_),
    .Y(_2194_));
 sky130_fd_sc_hd__nor2_1 _7106_ (.A(_2192_),
    .B(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__and2_1 _7107_ (.A(net11),
    .B(net40),
    .X(_2196_));
 sky130_fd_sc_hd__a21oi_1 _7108_ (.A1(_2192_),
    .A2(_2194_),
    .B1(_2196_),
    .Y(_2197_));
 sky130_fd_sc_hd__o31a_1 _7109_ (.A1(_2063_),
    .A2(_2195_),
    .A3(_2197_),
    .B1(_2065_),
    .X(_2198_));
 sky130_fd_sc_hd__xnor2_1 _7110_ (.A(_1906_),
    .B(_2050_),
    .Y(_2199_));
 sky130_fd_sc_hd__xnor2_2 _7111_ (.A(_2052_),
    .B(_2199_),
    .Y(_2201_));
 sky130_fd_sc_hd__nor2_1 _7112_ (.A(_2198_),
    .B(_2201_),
    .Y(_2202_));
 sky130_fd_sc_hd__nand2_1 _7113_ (.A(net14),
    .B(net40),
    .Y(_2203_));
 sky130_fd_sc_hd__a21oi_2 _7114_ (.A1(_2198_),
    .A2(_2201_),
    .B1(_2203_),
    .Y(_2204_));
 sky130_fd_sc_hd__o31ai_2 _7115_ (.A1(_2056_),
    .A2(_2202_),
    .A3(_2204_),
    .B1(_2059_),
    .Y(_2205_));
 sky130_fd_sc_hd__a31o_1 _7116_ (.A1(_1901_),
    .A2(_2051_),
    .A3(_2053_),
    .B1(_1902_),
    .X(_2206_));
 sky130_fd_sc_hd__nand2b_1 _7117_ (.A_N(_2206_),
    .B(_2205_),
    .Y(_2207_));
 sky130_fd_sc_hd__nor2_1 _7118_ (.A(_0099_),
    .B(_1727_),
    .Y(_2208_));
 sky130_fd_sc_hd__and2_1 _7119_ (.A(_2207_),
    .B(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__a21oi_1 _7120_ (.A1(net41),
    .A2(_1716_),
    .B1(_2209_),
    .Y(_2210_));
 sky130_fd_sc_hd__nand2_1 _7121_ (.A(net41),
    .B(_2209_),
    .Y(_2212_));
 sky130_fd_sc_hd__xnor2_1 _7122_ (.A(_3978_),
    .B(_2209_),
    .Y(_2213_));
 sky130_fd_sc_hd__xor2_1 _7123_ (.A(_2205_),
    .B(_2206_),
    .X(_2214_));
 sky130_fd_sc_hd__xnor2_1 _7124_ (.A(_2208_),
    .B(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__nand2_1 _7125_ (.A(net14),
    .B(net41),
    .Y(_2216_));
 sky130_fd_sc_hd__o22ai_2 _7126_ (.A1(_2056_),
    .A2(_2058_),
    .B1(_2202_),
    .B2(_2204_),
    .Y(_2217_));
 sky130_fd_sc_hd__or4_1 _7127_ (.A(_2056_),
    .B(_2058_),
    .C(_2202_),
    .D(_2204_),
    .X(_2218_));
 sky130_fd_sc_hd__and3_1 _7128_ (.A(_2216_),
    .B(_2217_),
    .C(_2218_),
    .X(_2219_));
 sky130_fd_sc_hd__nand3_1 _7129_ (.A(_2216_),
    .B(_2217_),
    .C(_2218_),
    .Y(_2220_));
 sky130_fd_sc_hd__a21oi_1 _7130_ (.A1(_2217_),
    .A2(_2218_),
    .B1(_2216_),
    .Y(_2221_));
 sky130_fd_sc_hd__and2_1 _7131_ (.A(net11),
    .B(net41),
    .X(_2223_));
 sky130_fd_sc_hd__o22ai_1 _7132_ (.A1(_2063_),
    .A2(_2064_),
    .B1(_2195_),
    .B2(_2197_),
    .Y(_2224_));
 sky130_fd_sc_hd__or4_1 _7133_ (.A(_2063_),
    .B(_2064_),
    .C(_2195_),
    .D(_2197_),
    .X(_2225_));
 sky130_fd_sc_hd__a21oi_1 _7134_ (.A1(_2224_),
    .A2(_2225_),
    .B1(_2223_),
    .Y(_2226_));
 sky130_fd_sc_hd__a21o_1 _7135_ (.A1(_2224_),
    .A2(_2225_),
    .B1(_2223_),
    .X(_2227_));
 sky130_fd_sc_hd__and3_1 _7136_ (.A(_2223_),
    .B(_2224_),
    .C(_2225_),
    .X(_2228_));
 sky130_fd_sc_hd__and2_1 _7137_ (.A(net9),
    .B(net41),
    .X(_2229_));
 sky130_fd_sc_hd__a2bb2o_1 _7138_ (.A1_N(_2070_),
    .A2_N(_2072_),
    .B1(_2188_),
    .B2(_2191_),
    .X(_2230_));
 sky130_fd_sc_hd__or4bb_1 _7139_ (.A(_2070_),
    .B(_2072_),
    .C_N(_2188_),
    .D_N(_2191_),
    .X(_2231_));
 sky130_fd_sc_hd__and3_1 _7140_ (.A(_2229_),
    .B(_2230_),
    .C(_2231_),
    .X(_2232_));
 sky130_fd_sc_hd__nand3_1 _7141_ (.A(_2229_),
    .B(_2230_),
    .C(_2231_),
    .Y(_2234_));
 sky130_fd_sc_hd__a21o_1 _7142_ (.A1(_2230_),
    .A2(_2231_),
    .B1(_2229_),
    .X(_2235_));
 sky130_fd_sc_hd__nand2_1 _7143_ (.A(net7),
    .B(net41),
    .Y(_2236_));
 sky130_fd_sc_hd__o211ai_2 _7144_ (.A1(_2076_),
    .A2(_2078_),
    .B1(_2182_),
    .C1(_2184_),
    .Y(_2237_));
 sky130_fd_sc_hd__a211o_1 _7145_ (.A1(_2182_),
    .A2(_2184_),
    .B1(_2076_),
    .C1(_2078_),
    .X(_2238_));
 sky130_fd_sc_hd__and3_1 _7146_ (.A(_2236_),
    .B(_2237_),
    .C(_2238_),
    .X(_2239_));
 sky130_fd_sc_hd__nand3_1 _7147_ (.A(_2236_),
    .B(_2237_),
    .C(_2238_),
    .Y(_2240_));
 sky130_fd_sc_hd__a21oi_1 _7148_ (.A1(_2237_),
    .A2(_2238_),
    .B1(_2236_),
    .Y(_2241_));
 sky130_fd_sc_hd__xor2_1 _7149_ (.A(_2179_),
    .B(_2181_),
    .X(_2242_));
 sky130_fd_sc_hd__xnor2_1 _7150_ (.A(_2183_),
    .B(_2242_),
    .Y(_2243_));
 sky130_fd_sc_hd__and2_1 _7151_ (.A(net5),
    .B(net41),
    .X(_2245_));
 sky130_fd_sc_hd__o211ai_2 _7152_ (.A1(_2083_),
    .A2(_2085_),
    .B1(_2175_),
    .C1(_2177_),
    .Y(_2246_));
 sky130_fd_sc_hd__a211o_1 _7153_ (.A1(_2175_),
    .A2(_2177_),
    .B1(_2083_),
    .C1(_2085_),
    .X(_2247_));
 sky130_fd_sc_hd__and3_1 _7154_ (.A(_2245_),
    .B(_2246_),
    .C(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__a21oi_1 _7155_ (.A1(_2246_),
    .A2(_2247_),
    .B1(_2245_),
    .Y(_2249_));
 sky130_fd_sc_hd__a21o_1 _7156_ (.A1(_2246_),
    .A2(_2247_),
    .B1(_2245_),
    .X(_2250_));
 sky130_fd_sc_hd__and2_1 _7157_ (.A(net3),
    .B(net41),
    .X(_2251_));
 sky130_fd_sc_hd__o211ai_1 _7158_ (.A1(_2089_),
    .A2(_2091_),
    .B1(_2169_),
    .C1(_2171_),
    .Y(_2252_));
 sky130_fd_sc_hd__a211o_1 _7159_ (.A1(_2169_),
    .A2(_2171_),
    .B1(_2089_),
    .C1(_2091_),
    .X(_2253_));
 sky130_fd_sc_hd__a21o_1 _7160_ (.A1(_2252_),
    .A2(_2253_),
    .B1(_2251_),
    .X(_2254_));
 sky130_fd_sc_hd__and3_1 _7161_ (.A(_2251_),
    .B(_2252_),
    .C(_2253_),
    .X(_2256_));
 sky130_fd_sc_hd__and2_1 _7162_ (.A(net32),
    .B(net41),
    .X(_2257_));
 sky130_fd_sc_hd__a22o_1 _7163_ (.A1(_2096_),
    .A2(_2098_),
    .B1(_2160_),
    .B2(_2163_),
    .X(_2258_));
 sky130_fd_sc_hd__nand4_1 _7164_ (.A(_2096_),
    .B(_2098_),
    .C(_2160_),
    .D(_2163_),
    .Y(_2259_));
 sky130_fd_sc_hd__a21oi_2 _7165_ (.A1(_2258_),
    .A2(_2259_),
    .B1(_2257_),
    .Y(_2260_));
 sky130_fd_sc_hd__and3_1 _7166_ (.A(_2257_),
    .B(_2258_),
    .C(_2259_),
    .X(_2261_));
 sky130_fd_sc_hd__and2_1 _7167_ (.A(net30),
    .B(net41),
    .X(_2262_));
 sky130_fd_sc_hd__xnor2_1 _7168_ (.A(_2100_),
    .B(_2102_),
    .Y(_2263_));
 sky130_fd_sc_hd__xnor2_2 _7169_ (.A(_2153_),
    .B(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hd__or2_1 _7170_ (.A(_2262_),
    .B(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__and2_1 _7171_ (.A(_2262_),
    .B(_2264_),
    .X(_2267_));
 sky130_fd_sc_hd__nand2_1 _7172_ (.A(net29),
    .B(net41),
    .Y(_2268_));
 sky130_fd_sc_hd__inv_2 _7173_ (.A(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__xnor2_1 _7174_ (.A(_2104_),
    .B(_2106_),
    .Y(_2270_));
 sky130_fd_sc_hd__xnor2_1 _7175_ (.A(_2151_),
    .B(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__or2_1 _7176_ (.A(_2269_),
    .B(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__and2_1 _7177_ (.A(net28),
    .B(net41),
    .X(_2273_));
 sky130_fd_sc_hd__o21bai_1 _7178_ (.A1(_2111_),
    .A2(_2113_),
    .B1_N(_2150_),
    .Y(_2274_));
 sky130_fd_sc_hd__or3b_1 _7179_ (.A(_2111_),
    .B(_2113_),
    .C_N(_2150_),
    .X(_2275_));
 sky130_fd_sc_hd__a21oi_1 _7180_ (.A1(_2274_),
    .A2(_2275_),
    .B1(_2273_),
    .Y(_2276_));
 sky130_fd_sc_hd__a21o_1 _7181_ (.A1(_2274_),
    .A2(_2275_),
    .B1(_2273_),
    .X(_2278_));
 sky130_fd_sc_hd__and3_1 _7182_ (.A(_2273_),
    .B(_2274_),
    .C(_2275_),
    .X(_2279_));
 sky130_fd_sc_hd__and2_1 _7183_ (.A(net27),
    .B(net41),
    .X(_2280_));
 sky130_fd_sc_hd__a22o_1 _7184_ (.A1(_2118_),
    .A2(_2120_),
    .B1(_2125_),
    .B2(_2149_),
    .X(_2281_));
 sky130_fd_sc_hd__nand4_1 _7185_ (.A(_2118_),
    .B(_2120_),
    .C(_2125_),
    .D(_2149_),
    .Y(_2282_));
 sky130_fd_sc_hd__a21oi_1 _7186_ (.A1(_2281_),
    .A2(_2282_),
    .B1(_2280_),
    .Y(_2283_));
 sky130_fd_sc_hd__a21o_1 _7187_ (.A1(_2281_),
    .A2(_2282_),
    .B1(_2280_),
    .X(_2284_));
 sky130_fd_sc_hd__and3_1 _7188_ (.A(_2280_),
    .B(_2281_),
    .C(_2282_),
    .X(_2285_));
 sky130_fd_sc_hd__nand2_1 _7189_ (.A(net26),
    .B(net41),
    .Y(_2286_));
 sky130_fd_sc_hd__xnor2_1 _7190_ (.A(_2121_),
    .B(_2124_),
    .Y(_2287_));
 sky130_fd_sc_hd__xnor2_1 _7191_ (.A(_2148_),
    .B(_2287_),
    .Y(_2289_));
 sky130_fd_sc_hd__nand2b_1 _7192_ (.A_N(_2289_),
    .B(_2286_),
    .Y(_2290_));
 sky130_fd_sc_hd__nand2_1 _7193_ (.A(net23),
    .B(net41),
    .Y(_2291_));
 sky130_fd_sc_hd__xor2_1 _7194_ (.A(_2126_),
    .B(_2128_),
    .X(_2292_));
 sky130_fd_sc_hd__xnor2_1 _7195_ (.A(_2146_),
    .B(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__nand2b_1 _7196_ (.A_N(_2293_),
    .B(_2291_),
    .Y(_2294_));
 sky130_fd_sc_hd__nand2_1 _7197_ (.A(net12),
    .B(net41),
    .Y(_2295_));
 sky130_fd_sc_hd__inv_2 _7198_ (.A(_2295_),
    .Y(_2296_));
 sky130_fd_sc_hd__xnor2_1 _7199_ (.A(_2130_),
    .B(_2132_),
    .Y(_2297_));
 sky130_fd_sc_hd__xnor2_1 _7200_ (.A(_2143_),
    .B(_2297_),
    .Y(_2298_));
 sky130_fd_sc_hd__and2_1 _7201_ (.A(_2296_),
    .B(_2298_),
    .X(_2300_));
 sky130_fd_sc_hd__nand2_1 _7202_ (.A(net1),
    .B(net41),
    .Y(_2301_));
 sky130_fd_sc_hd__or2_1 _7203_ (.A(_2138_),
    .B(_2141_),
    .X(_2302_));
 sky130_fd_sc_hd__a41o_1 _7204_ (.A1(_2135_),
    .A2(_2136_),
    .A3(_2137_),
    .A4(_2141_),
    .B1(_2301_),
    .X(_2303_));
 sky130_fd_sc_hd__a21oi_1 _7205_ (.A1(_2143_),
    .A2(_2302_),
    .B1(_2303_),
    .Y(_2304_));
 sky130_fd_sc_hd__o21a_1 _7206_ (.A1(_2296_),
    .A2(_2298_),
    .B1(_2304_),
    .X(_2305_));
 sky130_fd_sc_hd__nor2_1 _7207_ (.A(_2300_),
    .B(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__a311o_1 _7208_ (.A1(net23),
    .A2(net41),
    .A3(_2293_),
    .B1(_2300_),
    .C1(_2305_),
    .X(_2307_));
 sky130_fd_sc_hd__nand2_1 _7209_ (.A(_2294_),
    .B(_2307_),
    .Y(_2308_));
 sky130_fd_sc_hd__a32o_1 _7210_ (.A1(net26),
    .A2(net41),
    .A3(_2289_),
    .B1(_2294_),
    .B2(_2307_),
    .X(_2309_));
 sky130_fd_sc_hd__a31o_1 _7211_ (.A1(_2284_),
    .A2(_2290_),
    .A3(_2309_),
    .B1(_2285_),
    .X(_2311_));
 sky130_fd_sc_hd__a21oi_1 _7212_ (.A1(_2278_),
    .A2(_2311_),
    .B1(_2279_),
    .Y(_2312_));
 sky130_fd_sc_hd__a221o_1 _7213_ (.A1(_2269_),
    .A2(_2271_),
    .B1(_2278_),
    .B2(_2311_),
    .C1(_2279_),
    .X(_2313_));
 sky130_fd_sc_hd__nand2_1 _7214_ (.A(_2272_),
    .B(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__a22o_1 _7215_ (.A1(_2262_),
    .A2(_2264_),
    .B1(_2272_),
    .B2(_2313_),
    .X(_2315_));
 sky130_fd_sc_hd__o211a_1 _7216_ (.A1(_2262_),
    .A2(_2264_),
    .B1(_2272_),
    .C1(_2313_),
    .X(_2316_));
 sky130_fd_sc_hd__a21o_1 _7217_ (.A1(_2160_),
    .A2(_2161_),
    .B1(_2162_),
    .X(_2317_));
 sky130_fd_sc_hd__nand3_1 _7218_ (.A(_2160_),
    .B(_2161_),
    .C(_2162_),
    .Y(_2318_));
 sky130_fd_sc_hd__a211o_1 _7219_ (.A1(_2317_),
    .A2(_2318_),
    .B1(_2267_),
    .C1(_2316_),
    .X(_2319_));
 sky130_fd_sc_hd__o211ai_1 _7220_ (.A1(_2267_),
    .A2(_2316_),
    .B1(_2317_),
    .C1(_2318_),
    .Y(_2320_));
 sky130_fd_sc_hd__and2_1 _7221_ (.A(net31),
    .B(net41),
    .X(_2322_));
 sky130_fd_sc_hd__a41o_1 _7222_ (.A1(_2265_),
    .A2(_2315_),
    .A3(_2317_),
    .A4(_2318_),
    .B1(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__a21oi_2 _7223_ (.A1(_2319_),
    .A2(_2323_),
    .B1(_2261_),
    .Y(_2324_));
 sky130_fd_sc_hd__a21oi_2 _7224_ (.A1(_2168_),
    .A2(_2169_),
    .B1(_2170_),
    .Y(_2325_));
 sky130_fd_sc_hd__and3_1 _7225_ (.A(_2168_),
    .B(_2169_),
    .C(_2170_),
    .X(_2326_));
 sky130_fd_sc_hd__o22ai_4 _7226_ (.A1(_2260_),
    .A2(_2324_),
    .B1(_2325_),
    .B2(_2326_),
    .Y(_2327_));
 sky130_fd_sc_hd__or4_1 _7227_ (.A(_2260_),
    .B(_2324_),
    .C(_2325_),
    .D(_2326_),
    .X(_2328_));
 sky130_fd_sc_hd__and2_1 _7228_ (.A(net2),
    .B(net41),
    .X(_2329_));
 sky130_fd_sc_hd__nand2_1 _7229_ (.A(net2),
    .B(net41),
    .Y(_2330_));
 sky130_fd_sc_hd__o41ai_2 _7230_ (.A1(_2260_),
    .A2(_2324_),
    .A3(_2325_),
    .A4(_2326_),
    .B1(_2330_),
    .Y(_2331_));
 sky130_fd_sc_hd__a21o_1 _7231_ (.A1(_2327_),
    .A2(_2331_),
    .B1(_2256_),
    .X(_2333_));
 sky130_fd_sc_hd__a31o_1 _7232_ (.A1(_2254_),
    .A2(_2327_),
    .A3(_2331_),
    .B1(_2256_),
    .X(_2334_));
 sky130_fd_sc_hd__xor2_1 _7233_ (.A(_2172_),
    .B(_2174_),
    .X(_2335_));
 sky130_fd_sc_hd__xnor2_1 _7234_ (.A(_2176_),
    .B(_2335_),
    .Y(_2336_));
 sky130_fd_sc_hd__and2_1 _7235_ (.A(_2334_),
    .B(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__nand2_1 _7236_ (.A(net4),
    .B(net41),
    .Y(_2338_));
 sky130_fd_sc_hd__o211a_1 _7237_ (.A1(_2334_),
    .A2(_2336_),
    .B1(net4),
    .C1(net41),
    .X(_2339_));
 sky130_fd_sc_hd__o31a_1 _7238_ (.A1(_2248_),
    .A2(_2337_),
    .A3(_2339_),
    .B1(_2250_),
    .X(_2340_));
 sky130_fd_sc_hd__or2_1 _7239_ (.A(_2243_),
    .B(_2340_),
    .X(_2341_));
 sky130_fd_sc_hd__and2_1 _7240_ (.A(net6),
    .B(net41),
    .X(_2342_));
 sky130_fd_sc_hd__a21o_1 _7241_ (.A1(_2243_),
    .A2(_2340_),
    .B1(_2342_),
    .X(_2344_));
 sky130_fd_sc_hd__a31o_1 _7242_ (.A1(_2240_),
    .A2(_2341_),
    .A3(_2344_),
    .B1(_2241_),
    .X(_2345_));
 sky130_fd_sc_hd__xor2_1 _7243_ (.A(_2185_),
    .B(_2187_),
    .X(_2346_));
 sky130_fd_sc_hd__xnor2_1 _7244_ (.A(_2190_),
    .B(_2346_),
    .Y(_2347_));
 sky130_fd_sc_hd__or2_1 _7245_ (.A(_2345_),
    .B(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__nand2_1 _7246_ (.A(net8),
    .B(net41),
    .Y(_2349_));
 sky130_fd_sc_hd__a21bo_1 _7247_ (.A1(_2345_),
    .A2(_2347_),
    .B1_N(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__a31o_1 _7248_ (.A1(_2235_),
    .A2(_2348_),
    .A3(_2350_),
    .B1(_2232_),
    .X(_2351_));
 sky130_fd_sc_hd__xnor2_1 _7249_ (.A(_2192_),
    .B(_2194_),
    .Y(_2352_));
 sky130_fd_sc_hd__xnor2_1 _7250_ (.A(_2196_),
    .B(_2352_),
    .Y(_2353_));
 sky130_fd_sc_hd__or2_1 _7251_ (.A(_2351_),
    .B(_2353_),
    .X(_2355_));
 sky130_fd_sc_hd__and2_1 _7252_ (.A(net10),
    .B(net41),
    .X(_2356_));
 sky130_fd_sc_hd__a21o_1 _7253_ (.A1(_2351_),
    .A2(_2353_),
    .B1(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__a31o_1 _7254_ (.A1(_2227_),
    .A2(_2355_),
    .A3(_2357_),
    .B1(_2228_),
    .X(_2358_));
 sky130_fd_sc_hd__xor2_1 _7255_ (.A(_2198_),
    .B(_2201_),
    .X(_2359_));
 sky130_fd_sc_hd__xnor2_1 _7256_ (.A(_2203_),
    .B(_2359_),
    .Y(_2360_));
 sky130_fd_sc_hd__or2_1 _7257_ (.A(_2358_),
    .B(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__nand2_1 _7258_ (.A(net13),
    .B(net41),
    .Y(_2362_));
 sky130_fd_sc_hd__a21bo_1 _7259_ (.A1(_2358_),
    .A2(_2360_),
    .B1_N(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__a31o_1 _7260_ (.A1(_2220_),
    .A2(_2361_),
    .A3(_2363_),
    .B1(_2221_),
    .X(_2364_));
 sky130_fd_sc_hd__nor2_1 _7261_ (.A(_2215_),
    .B(_2364_),
    .Y(_2366_));
 sky130_fd_sc_hd__and2_1 _7262_ (.A(net15),
    .B(net41),
    .X(_2367_));
 sky130_fd_sc_hd__a21oi_1 _7263_ (.A1(_2215_),
    .A2(_2364_),
    .B1(_2367_),
    .Y(_2368_));
 sky130_fd_sc_hd__or3_1 _7264_ (.A(_2213_),
    .B(_2366_),
    .C(_2368_),
    .X(_2369_));
 sky130_fd_sc_hd__o21ai_1 _7265_ (.A1(_2366_),
    .A2(_2368_),
    .B1(_2213_),
    .Y(_2370_));
 sky130_fd_sc_hd__and3_1 _7266_ (.A(_3977_),
    .B(_2369_),
    .C(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__a21oi_1 _7267_ (.A1(_2369_),
    .A2(_2370_),
    .B1(_3977_),
    .Y(_2372_));
 sky130_fd_sc_hd__a21o_1 _7268_ (.A1(_2369_),
    .A2(_2370_),
    .B1(_3977_),
    .X(_2373_));
 sky130_fd_sc_hd__and2_1 _7269_ (.A(net13),
    .B(net42),
    .X(_2374_));
 sky130_fd_sc_hd__a2bb2o_1 _7270_ (.A1_N(_2219_),
    .A2_N(_2221_),
    .B1(_2361_),
    .B2(_2363_),
    .X(_2375_));
 sky130_fd_sc_hd__or4bb_1 _7271_ (.A(_2219_),
    .B(_2221_),
    .C_N(_2361_),
    .D_N(_2363_),
    .X(_2377_));
 sky130_fd_sc_hd__a21oi_1 _7272_ (.A1(_2375_),
    .A2(_2377_),
    .B1(_2374_),
    .Y(_2378_));
 sky130_fd_sc_hd__a21o_1 _7273_ (.A1(_2375_),
    .A2(_2377_),
    .B1(_2374_),
    .X(_2379_));
 sky130_fd_sc_hd__and3_1 _7274_ (.A(_2374_),
    .B(_2375_),
    .C(_2377_),
    .X(_2380_));
 sky130_fd_sc_hd__and2_1 _7275_ (.A(net10),
    .B(net42),
    .X(_2381_));
 sky130_fd_sc_hd__a2bb2o_1 _7276_ (.A1_N(_2226_),
    .A2_N(_2228_),
    .B1(_2355_),
    .B2(_2357_),
    .X(_2382_));
 sky130_fd_sc_hd__or4bb_1 _7277_ (.A(_2226_),
    .B(_2228_),
    .C_N(_2355_),
    .D_N(_2357_),
    .X(_2383_));
 sky130_fd_sc_hd__a21oi_1 _7278_ (.A1(_2382_),
    .A2(_2383_),
    .B1(_2381_),
    .Y(_2384_));
 sky130_fd_sc_hd__a21o_1 _7279_ (.A1(_2382_),
    .A2(_2383_),
    .B1(_2381_),
    .X(_2385_));
 sky130_fd_sc_hd__and3_1 _7280_ (.A(_2381_),
    .B(_2382_),
    .C(_2383_),
    .X(_2386_));
 sky130_fd_sc_hd__a22o_1 _7281_ (.A1(_2234_),
    .A2(_2235_),
    .B1(_2348_),
    .B2(_2350_),
    .X(_2388_));
 sky130_fd_sc_hd__nand4_1 _7282_ (.A(_2234_),
    .B(_2235_),
    .C(_2348_),
    .D(_2350_),
    .Y(_2389_));
 sky130_fd_sc_hd__a22oi_1 _7283_ (.A1(net8),
    .A2(net42),
    .B1(_2388_),
    .B2(_2389_),
    .Y(_2390_));
 sky130_fd_sc_hd__a22o_1 _7284_ (.A1(net8),
    .A2(net42),
    .B1(_2388_),
    .B2(_2389_),
    .X(_2391_));
 sky130_fd_sc_hd__and4_1 _7285_ (.A(net8),
    .B(net42),
    .C(_2388_),
    .D(_2389_),
    .X(_2392_));
 sky130_fd_sc_hd__and2_1 _7286_ (.A(net6),
    .B(net42),
    .X(_2393_));
 sky130_fd_sc_hd__a2bb2o_1 _7287_ (.A1_N(_2239_),
    .A2_N(_2241_),
    .B1(_2341_),
    .B2(_2344_),
    .X(_2394_));
 sky130_fd_sc_hd__or4bb_1 _7288_ (.A(_2239_),
    .B(_2241_),
    .C_N(_2341_),
    .D_N(_2344_),
    .X(_2395_));
 sky130_fd_sc_hd__a21oi_1 _7289_ (.A1(_2394_),
    .A2(_2395_),
    .B1(_2393_),
    .Y(_2396_));
 sky130_fd_sc_hd__a21o_1 _7290_ (.A1(_2394_),
    .A2(_2395_),
    .B1(_2393_),
    .X(_2397_));
 sky130_fd_sc_hd__and3_1 _7291_ (.A(_2393_),
    .B(_2394_),
    .C(_2395_),
    .X(_2399_));
 sky130_fd_sc_hd__nand2_1 _7292_ (.A(net4),
    .B(net42),
    .Y(_2400_));
 sky130_fd_sc_hd__o22ai_1 _7293_ (.A1(_2248_),
    .A2(_2249_),
    .B1(_2337_),
    .B2(_2339_),
    .Y(_2401_));
 sky130_fd_sc_hd__or4_1 _7294_ (.A(_2248_),
    .B(_2249_),
    .C(_2337_),
    .D(_2339_),
    .X(_2402_));
 sky130_fd_sc_hd__a21oi_1 _7295_ (.A1(_2401_),
    .A2(_2402_),
    .B1(_2400_),
    .Y(_2403_));
 sky130_fd_sc_hd__nand3_1 _7296_ (.A(_2400_),
    .B(_2401_),
    .C(_2402_),
    .Y(_2404_));
 sky130_fd_sc_hd__and2_1 _7297_ (.A(net2),
    .B(net42),
    .X(_2405_));
 sky130_fd_sc_hd__inv_2 _7298_ (.A(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__a21oi_1 _7299_ (.A1(_2327_),
    .A2(_2331_),
    .B1(_2254_),
    .Y(_2407_));
 sky130_fd_sc_hd__nand3_1 _7300_ (.A(_2256_),
    .B(_2327_),
    .C(_2331_),
    .Y(_2408_));
 sky130_fd_sc_hd__o211a_1 _7301_ (.A1(_2334_),
    .A2(_2407_),
    .B1(_2408_),
    .C1(_2406_),
    .X(_2410_));
 sky130_fd_sc_hd__a311o_1 _7302_ (.A1(_2254_),
    .A2(_2333_),
    .A3(_2408_),
    .B1(_2407_),
    .C1(_2406_),
    .X(_2411_));
 sky130_fd_sc_hd__and2_1 _7303_ (.A(net31),
    .B(net42),
    .X(_2412_));
 sky130_fd_sc_hd__or4bb_1 _7304_ (.A(_2260_),
    .B(_2261_),
    .C_N(_2319_),
    .D_N(_2323_),
    .X(_2413_));
 sky130_fd_sc_hd__a2bb2o_1 _7305_ (.A1_N(_2260_),
    .A2_N(_2261_),
    .B1(_2319_),
    .B2(_2323_),
    .X(_2414_));
 sky130_fd_sc_hd__a21oi_1 _7306_ (.A1(_2413_),
    .A2(_2414_),
    .B1(_2412_),
    .Y(_2415_));
 sky130_fd_sc_hd__a21o_1 _7307_ (.A1(_2413_),
    .A2(_2414_),
    .B1(_2412_),
    .X(_2416_));
 sky130_fd_sc_hd__and3_1 _7308_ (.A(_2412_),
    .B(_2413_),
    .C(_2414_),
    .X(_2417_));
 sky130_fd_sc_hd__and2_1 _7309_ (.A(net29),
    .B(net42),
    .X(_2418_));
 sky130_fd_sc_hd__xor2_1 _7310_ (.A(_2262_),
    .B(_2264_),
    .X(_2419_));
 sky130_fd_sc_hd__xnor2_1 _7311_ (.A(_2314_),
    .B(_2419_),
    .Y(_2421_));
 sky130_fd_sc_hd__or2_1 _7312_ (.A(_2418_),
    .B(_2421_),
    .X(_2422_));
 sky130_fd_sc_hd__nand2_1 _7313_ (.A(net28),
    .B(net42),
    .Y(_2423_));
 sky130_fd_sc_hd__inv_2 _7314_ (.A(_2423_),
    .Y(_2424_));
 sky130_fd_sc_hd__xnor2_1 _7315_ (.A(_2268_),
    .B(_2271_),
    .Y(_2425_));
 sky130_fd_sc_hd__xnor2_1 _7316_ (.A(_2312_),
    .B(_2425_),
    .Y(_2426_));
 sky130_fd_sc_hd__or2_1 _7317_ (.A(_2424_),
    .B(_2426_),
    .X(_2427_));
 sky130_fd_sc_hd__nand2_1 _7318_ (.A(net27),
    .B(net42),
    .Y(_2428_));
 sky130_fd_sc_hd__o21ai_1 _7319_ (.A1(_2276_),
    .A2(_2279_),
    .B1(_2311_),
    .Y(_2429_));
 sky130_fd_sc_hd__or3_1 _7320_ (.A(_2276_),
    .B(_2279_),
    .C(_2311_),
    .X(_2430_));
 sky130_fd_sc_hd__and3_1 _7321_ (.A(_2428_),
    .B(_2429_),
    .C(_2430_),
    .X(_2432_));
 sky130_fd_sc_hd__nand3_1 _7322_ (.A(_2428_),
    .B(_2429_),
    .C(_2430_),
    .Y(_2433_));
 sky130_fd_sc_hd__a21oi_1 _7323_ (.A1(_2429_),
    .A2(_2430_),
    .B1(_2428_),
    .Y(_2434_));
 sky130_fd_sc_hd__and2_1 _7324_ (.A(net26),
    .B(net42),
    .X(_2435_));
 sky130_fd_sc_hd__or4bb_1 _7325_ (.A(_2283_),
    .B(_2285_),
    .C_N(_2290_),
    .D_N(_2309_),
    .X(_2436_));
 sky130_fd_sc_hd__a2bb2o_1 _7326_ (.A1_N(_2283_),
    .A2_N(_2285_),
    .B1(_2290_),
    .B2(_2309_),
    .X(_2437_));
 sky130_fd_sc_hd__and3_1 _7327_ (.A(_2435_),
    .B(_2436_),
    .C(_2437_),
    .X(_2438_));
 sky130_fd_sc_hd__a21oi_1 _7328_ (.A1(_2436_),
    .A2(_2437_),
    .B1(_2435_),
    .Y(_2439_));
 sky130_fd_sc_hd__a21o_1 _7329_ (.A1(_2436_),
    .A2(_2437_),
    .B1(_2435_),
    .X(_2440_));
 sky130_fd_sc_hd__nand2_1 _7330_ (.A(net23),
    .B(net42),
    .Y(_2441_));
 sky130_fd_sc_hd__xnor2_1 _7331_ (.A(_2286_),
    .B(_2289_),
    .Y(_2443_));
 sky130_fd_sc_hd__xnor2_1 _7332_ (.A(_2308_),
    .B(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__a21o_1 _7333_ (.A1(net23),
    .A2(net42),
    .B1(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__and2_1 _7334_ (.A(net12),
    .B(net42),
    .X(_2446_));
 sky130_fd_sc_hd__xnor2_1 _7335_ (.A(_2291_),
    .B(_2293_),
    .Y(_2447_));
 sky130_fd_sc_hd__xnor2_1 _7336_ (.A(_2306_),
    .B(_2447_),
    .Y(_2448_));
 sky130_fd_sc_hd__and2_1 _7337_ (.A(_2446_),
    .B(_2448_),
    .X(_2449_));
 sky130_fd_sc_hd__xnor2_1 _7338_ (.A(_2295_),
    .B(_2298_),
    .Y(_2450_));
 sky130_fd_sc_hd__or2_1 _7339_ (.A(_2304_),
    .B(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__nand2_1 _7340_ (.A(_2304_),
    .B(_2450_),
    .Y(_2452_));
 sky130_fd_sc_hd__and4_1 _7341_ (.A(net1),
    .B(net42),
    .C(_2451_),
    .D(_2452_),
    .X(_2454_));
 sky130_fd_sc_hd__o21a_1 _7342_ (.A1(_2446_),
    .A2(_2448_),
    .B1(_2454_),
    .X(_2455_));
 sky130_fd_sc_hd__or2_1 _7343_ (.A(_2449_),
    .B(_2455_),
    .X(_2456_));
 sky130_fd_sc_hd__a311o_1 _7344_ (.A1(net23),
    .A2(net42),
    .A3(_2444_),
    .B1(_2449_),
    .C1(_2455_),
    .X(_2457_));
 sky130_fd_sc_hd__a31o_1 _7345_ (.A1(_2440_),
    .A2(_2445_),
    .A3(_2457_),
    .B1(_2438_),
    .X(_2458_));
 sky130_fd_sc_hd__a21oi_1 _7346_ (.A1(_2433_),
    .A2(_2458_),
    .B1(_2434_),
    .Y(_2459_));
 sky130_fd_sc_hd__a221o_1 _7347_ (.A1(_2424_),
    .A2(_2426_),
    .B1(_2433_),
    .B2(_2458_),
    .C1(_2434_),
    .X(_2460_));
 sky130_fd_sc_hd__nand2_1 _7348_ (.A(_2427_),
    .B(_2460_),
    .Y(_2461_));
 sky130_fd_sc_hd__a22o_1 _7349_ (.A1(_2418_),
    .A2(_2421_),
    .B1(_2427_),
    .B2(_2460_),
    .X(_2462_));
 sky130_fd_sc_hd__a21o_1 _7350_ (.A1(_2319_),
    .A2(_2320_),
    .B1(_2322_),
    .X(_2463_));
 sky130_fd_sc_hd__nand4_1 _7351_ (.A(net31),
    .B(net41),
    .C(_2319_),
    .D(_2320_),
    .Y(_2465_));
 sky130_fd_sc_hd__a22o_1 _7352_ (.A1(_2422_),
    .A2(_2462_),
    .B1(_2463_),
    .B2(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__nand4_1 _7353_ (.A(_2422_),
    .B(_2462_),
    .C(_2463_),
    .D(_2465_),
    .Y(_2467_));
 sky130_fd_sc_hd__nand2_1 _7354_ (.A(net30),
    .B(net42),
    .Y(_2468_));
 sky130_fd_sc_hd__inv_2 _7355_ (.A(_2468_),
    .Y(_2469_));
 sky130_fd_sc_hd__a41o_1 _7356_ (.A1(_2422_),
    .A2(_2462_),
    .A3(_2463_),
    .A4(_2465_),
    .B1(_2469_),
    .X(_2470_));
 sky130_fd_sc_hd__and2_1 _7357_ (.A(_2466_),
    .B(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__a31o_1 _7358_ (.A1(_2416_),
    .A2(_2466_),
    .A3(_2470_),
    .B1(_2417_),
    .X(_2472_));
 sky130_fd_sc_hd__a21o_1 _7359_ (.A1(_2327_),
    .A2(_2328_),
    .B1(_2329_),
    .X(_2473_));
 sky130_fd_sc_hd__nand3_1 _7360_ (.A(_2327_),
    .B(_2328_),
    .C(_2329_),
    .Y(_2474_));
 sky130_fd_sc_hd__a21oi_1 _7361_ (.A1(_2473_),
    .A2(_2474_),
    .B1(_2472_),
    .Y(_2476_));
 sky130_fd_sc_hd__and3_1 _7362_ (.A(_2472_),
    .B(_2473_),
    .C(_2474_),
    .X(_2477_));
 sky130_fd_sc_hd__and2_1 _7363_ (.A(net32),
    .B(net42),
    .X(_2478_));
 sky130_fd_sc_hd__a31oi_1 _7364_ (.A1(_2472_),
    .A2(_2473_),
    .A3(_2474_),
    .B1(_2478_),
    .Y(_2479_));
 sky130_fd_sc_hd__or2_1 _7365_ (.A(_2476_),
    .B(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__o31ai_1 _7366_ (.A1(_2410_),
    .A2(_2476_),
    .A3(_2479_),
    .B1(_2411_),
    .Y(_2481_));
 sky130_fd_sc_hd__xor2_1 _7367_ (.A(_2334_),
    .B(_2336_),
    .X(_2482_));
 sky130_fd_sc_hd__xnor2_1 _7368_ (.A(_2338_),
    .B(_2482_),
    .Y(_2483_));
 sky130_fd_sc_hd__or2_1 _7369_ (.A(_2481_),
    .B(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__nand2_1 _7370_ (.A(_2481_),
    .B(_2483_),
    .Y(_2485_));
 sky130_fd_sc_hd__and2_1 _7371_ (.A(net3),
    .B(net42),
    .X(_2487_));
 sky130_fd_sc_hd__a21o_1 _7372_ (.A1(_2481_),
    .A2(_2483_),
    .B1(_2487_),
    .X(_2488_));
 sky130_fd_sc_hd__nand2_1 _7373_ (.A(_2484_),
    .B(_2488_),
    .Y(_2489_));
 sky130_fd_sc_hd__a31o_1 _7374_ (.A1(_2404_),
    .A2(_2484_),
    .A3(_2488_),
    .B1(_2403_),
    .X(_2490_));
 sky130_fd_sc_hd__xnor2_1 _7375_ (.A(_2243_),
    .B(_2340_),
    .Y(_2491_));
 sky130_fd_sc_hd__xnor2_1 _7376_ (.A(_2342_),
    .B(_2491_),
    .Y(_2492_));
 sky130_fd_sc_hd__or2_1 _7377_ (.A(_2490_),
    .B(_2492_),
    .X(_2493_));
 sky130_fd_sc_hd__nand2_1 _7378_ (.A(net5),
    .B(net42),
    .Y(_2494_));
 sky130_fd_sc_hd__inv_2 _7379_ (.A(_2494_),
    .Y(_2495_));
 sky130_fd_sc_hd__a21o_1 _7380_ (.A1(_2490_),
    .A2(_2492_),
    .B1(_2495_),
    .X(_2496_));
 sky130_fd_sc_hd__a31o_1 _7381_ (.A1(_2397_),
    .A2(_2493_),
    .A3(_2496_),
    .B1(_2399_),
    .X(_2498_));
 sky130_fd_sc_hd__xor2_1 _7382_ (.A(_2345_),
    .B(_2347_),
    .X(_2499_));
 sky130_fd_sc_hd__xnor2_1 _7383_ (.A(_2349_),
    .B(_2499_),
    .Y(_2500_));
 sky130_fd_sc_hd__or2_1 _7384_ (.A(_2498_),
    .B(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__and2_1 _7385_ (.A(net7),
    .B(net42),
    .X(_2502_));
 sky130_fd_sc_hd__a21o_1 _7386_ (.A1(_2498_),
    .A2(_2500_),
    .B1(_2502_),
    .X(_2503_));
 sky130_fd_sc_hd__a31o_1 _7387_ (.A1(_2391_),
    .A2(_2501_),
    .A3(_2503_),
    .B1(_2392_),
    .X(_2504_));
 sky130_fd_sc_hd__xnor2_1 _7388_ (.A(_2351_),
    .B(_2353_),
    .Y(_2505_));
 sky130_fd_sc_hd__xnor2_1 _7389_ (.A(_2356_),
    .B(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__or2_1 _7390_ (.A(_2504_),
    .B(_2506_),
    .X(_2507_));
 sky130_fd_sc_hd__nand2_1 _7391_ (.A(net9),
    .B(net42),
    .Y(_2509_));
 sky130_fd_sc_hd__a21bo_1 _7392_ (.A1(_2504_),
    .A2(_2506_),
    .B1_N(_2509_),
    .X(_2510_));
 sky130_fd_sc_hd__a31o_1 _7393_ (.A1(_2385_),
    .A2(_2507_),
    .A3(_2510_),
    .B1(_2386_),
    .X(_2511_));
 sky130_fd_sc_hd__xor2_1 _7394_ (.A(_2358_),
    .B(_2360_),
    .X(_2512_));
 sky130_fd_sc_hd__xnor2_1 _7395_ (.A(_2362_),
    .B(_2512_),
    .Y(_2513_));
 sky130_fd_sc_hd__or2_1 _7396_ (.A(_2511_),
    .B(_2513_),
    .X(_2514_));
 sky130_fd_sc_hd__nand2_1 _7397_ (.A(net11),
    .B(net42),
    .Y(_2515_));
 sky130_fd_sc_hd__a21bo_1 _7398_ (.A1(_2511_),
    .A2(_2513_),
    .B1_N(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__a31o_1 _7399_ (.A1(_2379_),
    .A2(_2514_),
    .A3(_2516_),
    .B1(_2380_),
    .X(_2517_));
 sky130_fd_sc_hd__xnor2_1 _7400_ (.A(_2215_),
    .B(_2364_),
    .Y(_2518_));
 sky130_fd_sc_hd__xnor2_2 _7401_ (.A(_2367_),
    .B(_2518_),
    .Y(_2520_));
 sky130_fd_sc_hd__nor2_1 _7402_ (.A(_2517_),
    .B(_2520_),
    .Y(_2521_));
 sky130_fd_sc_hd__and2_1 _7403_ (.A(net14),
    .B(net42),
    .X(_2522_));
 sky130_fd_sc_hd__a21oi_1 _7404_ (.A1(_2517_),
    .A2(_2520_),
    .B1(_2522_),
    .Y(_2523_));
 sky130_fd_sc_hd__o31a_1 _7405_ (.A1(_2371_),
    .A2(_2521_),
    .A3(_2523_),
    .B1(_2373_),
    .X(_2524_));
 sky130_fd_sc_hd__o31a_1 _7406_ (.A1(_2210_),
    .A2(_2366_),
    .A3(_2368_),
    .B1(_2212_),
    .X(_2525_));
 sky130_fd_sc_hd__a21oi_1 _7407_ (.A1(_2524_),
    .A2(_2525_),
    .B1(_3976_),
    .Y(_2526_));
 sky130_fd_sc_hd__a21o_1 _7408_ (.A1(net43),
    .A2(_1716_),
    .B1(_2526_),
    .X(_2527_));
 sky130_fd_sc_hd__a21boi_1 _7409_ (.A1(net43),
    .A2(_2526_),
    .B1_N(_2527_),
    .Y(_2528_));
 sky130_fd_sc_hd__and2_1 _7410_ (.A(net14),
    .B(net43),
    .X(_2529_));
 sky130_fd_sc_hd__o22ai_2 _7411_ (.A1(_2371_),
    .A2(_2372_),
    .B1(_2521_),
    .B2(_2523_),
    .Y(_2531_));
 sky130_fd_sc_hd__or4_1 _7412_ (.A(_2371_),
    .B(_2372_),
    .C(_2521_),
    .D(_2523_),
    .X(_2532_));
 sky130_fd_sc_hd__a21o_1 _7413_ (.A1(_2531_),
    .A2(_2532_),
    .B1(_2529_),
    .X(_2533_));
 sky130_fd_sc_hd__and3_1 _7414_ (.A(_2529_),
    .B(_2531_),
    .C(_2532_),
    .X(_2534_));
 sky130_fd_sc_hd__nand3_1 _7415_ (.A(_2529_),
    .B(_2531_),
    .C(_2532_),
    .Y(_2535_));
 sky130_fd_sc_hd__nand2_1 _7416_ (.A(net11),
    .B(net43),
    .Y(_2536_));
 sky130_fd_sc_hd__o211ai_2 _7417_ (.A1(_2378_),
    .A2(_2380_),
    .B1(_2514_),
    .C1(_2516_),
    .Y(_2537_));
 sky130_fd_sc_hd__a211o_1 _7418_ (.A1(_2514_),
    .A2(_2516_),
    .B1(_2378_),
    .C1(_2380_),
    .X(_2538_));
 sky130_fd_sc_hd__and3_1 _7419_ (.A(_2536_),
    .B(_2537_),
    .C(_2538_),
    .X(_2539_));
 sky130_fd_sc_hd__a21oi_1 _7420_ (.A1(_2537_),
    .A2(_2538_),
    .B1(_2536_),
    .Y(_2540_));
 sky130_fd_sc_hd__a21o_1 _7421_ (.A1(_2537_),
    .A2(_2538_),
    .B1(_2536_),
    .X(_2542_));
 sky130_fd_sc_hd__xor2_1 _7422_ (.A(_2511_),
    .B(_2513_),
    .X(_2543_));
 sky130_fd_sc_hd__xnor2_2 _7423_ (.A(_2515_),
    .B(_2543_),
    .Y(_2544_));
 sky130_fd_sc_hd__and2_1 _7424_ (.A(net9),
    .B(net43),
    .X(_2545_));
 sky130_fd_sc_hd__a2bb2o_1 _7425_ (.A1_N(_2384_),
    .A2_N(_2386_),
    .B1(_2507_),
    .B2(_2510_),
    .X(_2546_));
 sky130_fd_sc_hd__or4bb_1 _7426_ (.A(_2384_),
    .B(_2386_),
    .C_N(_2507_),
    .D_N(_2510_),
    .X(_2547_));
 sky130_fd_sc_hd__a21oi_1 _7427_ (.A1(_2546_),
    .A2(_2547_),
    .B1(_2545_),
    .Y(_2548_));
 sky130_fd_sc_hd__a21o_1 _7428_ (.A1(_2546_),
    .A2(_2547_),
    .B1(_2545_),
    .X(_2549_));
 sky130_fd_sc_hd__and3_1 _7429_ (.A(_2545_),
    .B(_2546_),
    .C(_2547_),
    .X(_2550_));
 sky130_fd_sc_hd__xor2_1 _7430_ (.A(_2504_),
    .B(_2506_),
    .X(_2551_));
 sky130_fd_sc_hd__xnor2_1 _7431_ (.A(_2509_),
    .B(_2551_),
    .Y(_2553_));
 sky130_fd_sc_hd__and2_1 _7432_ (.A(net7),
    .B(net43),
    .X(_2554_));
 sky130_fd_sc_hd__a2bb2o_1 _7433_ (.A1_N(_2390_),
    .A2_N(_2392_),
    .B1(_2501_),
    .B2(_2503_),
    .X(_2555_));
 sky130_fd_sc_hd__or4bb_1 _7434_ (.A(_2390_),
    .B(_2392_),
    .C_N(_2501_),
    .D_N(_2503_),
    .X(_2556_));
 sky130_fd_sc_hd__and3_1 _7435_ (.A(_2554_),
    .B(_2555_),
    .C(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__a21o_1 _7436_ (.A1(_2555_),
    .A2(_2556_),
    .B1(_2554_),
    .X(_2558_));
 sky130_fd_sc_hd__nand2_2 _7437_ (.A(net5),
    .B(net43),
    .Y(_2559_));
 sky130_fd_sc_hd__o211a_1 _7438_ (.A1(_2396_),
    .A2(_2399_),
    .B1(_2493_),
    .C1(_2496_),
    .X(_2560_));
 sky130_fd_sc_hd__a211o_1 _7439_ (.A1(_2493_),
    .A2(_2496_),
    .B1(_2396_),
    .C1(_2399_),
    .X(_2561_));
 sky130_fd_sc_hd__and2b_1 _7440_ (.A_N(_2560_),
    .B(_2561_),
    .X(_2562_));
 sky130_fd_sc_hd__nor2_1 _7441_ (.A(_2559_),
    .B(_2562_),
    .Y(_2564_));
 sky130_fd_sc_hd__nand2_1 _7442_ (.A(net3),
    .B(net43),
    .Y(_2565_));
 sky130_fd_sc_hd__and2b_1 _7443_ (.A_N(_2403_),
    .B(_2404_),
    .X(_2566_));
 sky130_fd_sc_hd__xnor2_1 _7444_ (.A(_2489_),
    .B(_2566_),
    .Y(_2567_));
 sky130_fd_sc_hd__a21oi_1 _7445_ (.A1(net3),
    .A2(net43),
    .B1(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__nand2b_1 _7446_ (.A_N(_2565_),
    .B(_2567_),
    .Y(_2569_));
 sky130_fd_sc_hd__nand2_1 _7447_ (.A(net32),
    .B(net43),
    .Y(_2570_));
 sky130_fd_sc_hd__and2b_1 _7448_ (.A_N(_2410_),
    .B(_2411_),
    .X(_2571_));
 sky130_fd_sc_hd__xor2_1 _7449_ (.A(_2480_),
    .B(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__nand2_1 _7450_ (.A(_2570_),
    .B(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__nor2_1 _7451_ (.A(_2570_),
    .B(_2572_),
    .Y(_2575_));
 sky130_fd_sc_hd__nand2_1 _7452_ (.A(net30),
    .B(net43),
    .Y(_2576_));
 sky130_fd_sc_hd__or2_1 _7453_ (.A(_2415_),
    .B(_2417_),
    .X(_2577_));
 sky130_fd_sc_hd__xnor2_1 _7454_ (.A(_2471_),
    .B(_2577_),
    .Y(_2578_));
 sky130_fd_sc_hd__a21o_1 _7455_ (.A1(net30),
    .A2(net43),
    .B1(_2578_),
    .X(_2579_));
 sky130_fd_sc_hd__and3_1 _7456_ (.A(net30),
    .B(net43),
    .C(_2578_),
    .X(_2580_));
 sky130_fd_sc_hd__nand2_1 _7457_ (.A(net28),
    .B(net43),
    .Y(_2581_));
 sky130_fd_sc_hd__xor2_1 _7458_ (.A(_2418_),
    .B(_2421_),
    .X(_2582_));
 sky130_fd_sc_hd__xnor2_1 _7459_ (.A(_2461_),
    .B(_2582_),
    .Y(_2583_));
 sky130_fd_sc_hd__and3_1 _7460_ (.A(net28),
    .B(net43),
    .C(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__nand2b_1 _7461_ (.A_N(_2583_),
    .B(_2581_),
    .Y(_2586_));
 sky130_fd_sc_hd__and2_1 _7462_ (.A(net27),
    .B(net43),
    .X(_2587_));
 sky130_fd_sc_hd__xnor2_1 _7463_ (.A(_2423_),
    .B(_2426_),
    .Y(_2588_));
 sky130_fd_sc_hd__xnor2_1 _7464_ (.A(_2459_),
    .B(_2588_),
    .Y(_2589_));
 sky130_fd_sc_hd__nor2_1 _7465_ (.A(_2587_),
    .B(_2589_),
    .Y(_2590_));
 sky130_fd_sc_hd__nand2_1 _7466_ (.A(_2587_),
    .B(_2589_),
    .Y(_2591_));
 sky130_fd_sc_hd__and2_1 _7467_ (.A(net26),
    .B(net43),
    .X(_2592_));
 sky130_fd_sc_hd__o21bai_1 _7468_ (.A1(_2432_),
    .A2(_2434_),
    .B1_N(_2458_),
    .Y(_2593_));
 sky130_fd_sc_hd__or3b_1 _7469_ (.A(_2432_),
    .B(_2434_),
    .C_N(_2458_),
    .X(_2594_));
 sky130_fd_sc_hd__a21oi_1 _7470_ (.A1(_2593_),
    .A2(_2594_),
    .B1(_2592_),
    .Y(_2595_));
 sky130_fd_sc_hd__and3_1 _7471_ (.A(_2592_),
    .B(_2593_),
    .C(_2594_),
    .X(_2597_));
 sky130_fd_sc_hd__nand3_1 _7472_ (.A(_2592_),
    .B(_2593_),
    .C(_2594_),
    .Y(_2598_));
 sky130_fd_sc_hd__nand2_1 _7473_ (.A(net23),
    .B(net43),
    .Y(_2599_));
 sky130_fd_sc_hd__o211ai_1 _7474_ (.A1(_2438_),
    .A2(_2439_),
    .B1(_2445_),
    .C1(_2457_),
    .Y(_2600_));
 sky130_fd_sc_hd__a211o_1 _7475_ (.A1(_2445_),
    .A2(_2457_),
    .B1(_2438_),
    .C1(_2439_),
    .X(_2601_));
 sky130_fd_sc_hd__and3_1 _7476_ (.A(_2599_),
    .B(_2600_),
    .C(_2601_),
    .X(_2602_));
 sky130_fd_sc_hd__a21oi_2 _7477_ (.A1(_2600_),
    .A2(_2601_),
    .B1(_2599_),
    .Y(_2603_));
 sky130_fd_sc_hd__nand2_1 _7478_ (.A(net12),
    .B(net43),
    .Y(_2604_));
 sky130_fd_sc_hd__xnor2_1 _7479_ (.A(_2441_),
    .B(_2444_),
    .Y(_2605_));
 sky130_fd_sc_hd__xnor2_1 _7480_ (.A(_2456_),
    .B(_2605_),
    .Y(_2606_));
 sky130_fd_sc_hd__or2_2 _7481_ (.A(_2604_),
    .B(_2606_),
    .X(_2608_));
 sky130_fd_sc_hd__nand2_1 _7482_ (.A(_2604_),
    .B(_2606_),
    .Y(_2609_));
 sky130_fd_sc_hd__xor2_1 _7483_ (.A(_2446_),
    .B(_2448_),
    .X(_2610_));
 sky130_fd_sc_hd__nand2_1 _7484_ (.A(net1),
    .B(net43),
    .Y(_2611_));
 sky130_fd_sc_hd__a21oi_1 _7485_ (.A1(_2454_),
    .A2(_2610_),
    .B1(_2611_),
    .Y(_2612_));
 sky130_fd_sc_hd__o21ai_1 _7486_ (.A1(_2454_),
    .A2(_2610_),
    .B1(_2612_),
    .Y(_2613_));
 sky130_fd_sc_hd__a21o_1 _7487_ (.A1(_2604_),
    .A2(_2606_),
    .B1(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__and3b_1 _7488_ (.A_N(_2603_),
    .B(_2608_),
    .C(_2614_),
    .X(_2615_));
 sky130_fd_sc_hd__a21oi_1 _7489_ (.A1(_2608_),
    .A2(_2614_),
    .B1(_2602_),
    .Y(_2616_));
 sky130_fd_sc_hd__o31a_1 _7490_ (.A1(_2595_),
    .A2(_2602_),
    .A3(_2615_),
    .B1(_2598_),
    .X(_2617_));
 sky130_fd_sc_hd__o21ai_1 _7491_ (.A1(_2590_),
    .A2(_2617_),
    .B1(_2591_),
    .Y(_2619_));
 sky130_fd_sc_hd__a21o_1 _7492_ (.A1(_2586_),
    .A2(_2619_),
    .B1(_2584_),
    .X(_2620_));
 sky130_fd_sc_hd__nand2_1 _7493_ (.A(_2466_),
    .B(_2467_),
    .Y(_2621_));
 sky130_fd_sc_hd__xnor2_1 _7494_ (.A(_2469_),
    .B(_2621_),
    .Y(_2622_));
 sky130_fd_sc_hd__or2_1 _7495_ (.A(_2620_),
    .B(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__nand2_1 _7496_ (.A(net29),
    .B(net43),
    .Y(_2624_));
 sky130_fd_sc_hd__a21bo_1 _7497_ (.A1(_2620_),
    .A2(_2622_),
    .B1_N(_2624_),
    .X(_2625_));
 sky130_fd_sc_hd__a31o_1 _7498_ (.A1(_2579_),
    .A2(_2623_),
    .A3(_2625_),
    .B1(_2580_),
    .X(_2626_));
 sky130_fd_sc_hd__or2_1 _7499_ (.A(_2476_),
    .B(_2477_),
    .X(_2627_));
 sky130_fd_sc_hd__xnor2_2 _7500_ (.A(_2478_),
    .B(_2627_),
    .Y(_2628_));
 sky130_fd_sc_hd__or2_1 _7501_ (.A(_2626_),
    .B(_2628_),
    .X(_2630_));
 sky130_fd_sc_hd__nand2_1 _7502_ (.A(_2626_),
    .B(_2628_),
    .Y(_2631_));
 sky130_fd_sc_hd__and2_1 _7503_ (.A(net31),
    .B(net43),
    .X(_2632_));
 sky130_fd_sc_hd__a21o_1 _7504_ (.A1(_2626_),
    .A2(_2628_),
    .B1(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__o21ai_1 _7505_ (.A1(_2626_),
    .A2(_2628_),
    .B1(_2632_),
    .Y(_2634_));
 sky130_fd_sc_hd__a31o_1 _7506_ (.A1(_2573_),
    .A2(_2630_),
    .A3(_2633_),
    .B1(_2575_),
    .X(_2635_));
 sky130_fd_sc_hd__nand2_1 _7507_ (.A(_2484_),
    .B(_2485_),
    .Y(_2636_));
 sky130_fd_sc_hd__xnor2_2 _7508_ (.A(_2487_),
    .B(_2636_),
    .Y(_2637_));
 sky130_fd_sc_hd__nor2_1 _7509_ (.A(_2635_),
    .B(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__nand2_1 _7510_ (.A(_2635_),
    .B(_2637_),
    .Y(_2639_));
 sky130_fd_sc_hd__and2_1 _7511_ (.A(net2),
    .B(net43),
    .X(_2641_));
 sky130_fd_sc_hd__a21oi_1 _7512_ (.A1(_2635_),
    .A2(_2637_),
    .B1(_2641_),
    .Y(_2642_));
 sky130_fd_sc_hd__o211ai_1 _7513_ (.A1(_2635_),
    .A2(_2637_),
    .B1(net2),
    .C1(net43),
    .Y(_2643_));
 sky130_fd_sc_hd__xor2_1 _7514_ (.A(_2490_),
    .B(_2492_),
    .X(_2644_));
 sky130_fd_sc_hd__xnor2_1 _7515_ (.A(_2495_),
    .B(_2644_),
    .Y(_2645_));
 sky130_fd_sc_hd__o311a_1 _7516_ (.A1(_2568_),
    .A2(_2638_),
    .A3(_2642_),
    .B1(_2645_),
    .C1(_2569_),
    .X(_2646_));
 sky130_fd_sc_hd__a311o_1 _7517_ (.A1(_2569_),
    .A2(_2639_),
    .A3(_2643_),
    .B1(_2645_),
    .C1(_2568_),
    .X(_2647_));
 sky130_fd_sc_hd__nand2_2 _7518_ (.A(net4),
    .B(net43),
    .Y(_2648_));
 sky130_fd_sc_hd__a21oi_1 _7519_ (.A1(_2647_),
    .A2(_2648_),
    .B1(_2646_),
    .Y(_2649_));
 sky130_fd_sc_hd__a221oi_4 _7520_ (.A1(_2559_),
    .A2(_2562_),
    .B1(_2647_),
    .B2(_2648_),
    .C1(_2646_),
    .Y(_2650_));
 sky130_fd_sc_hd__xnor2_1 _7521_ (.A(_2498_),
    .B(_2500_),
    .Y(_2652_));
 sky130_fd_sc_hd__xnor2_1 _7522_ (.A(_2502_),
    .B(_2652_),
    .Y(_2653_));
 sky130_fd_sc_hd__nor3_1 _7523_ (.A(_2564_),
    .B(_2650_),
    .C(_2653_),
    .Y(_2654_));
 sky130_fd_sc_hd__o21a_1 _7524_ (.A1(_2564_),
    .A2(_2650_),
    .B1(_2653_),
    .X(_2655_));
 sky130_fd_sc_hd__nand2_1 _7525_ (.A(net6),
    .B(net43),
    .Y(_2656_));
 sky130_fd_sc_hd__o311a_1 _7526_ (.A1(_2564_),
    .A2(_2650_),
    .A3(_2653_),
    .B1(net43),
    .C1(net6),
    .X(_2657_));
 sky130_fd_sc_hd__nor2_1 _7527_ (.A(_2655_),
    .B(_2657_),
    .Y(_2658_));
 sky130_fd_sc_hd__o31a_1 _7528_ (.A1(_2557_),
    .A2(_2655_),
    .A3(_2657_),
    .B1(_2558_),
    .X(_2659_));
 sky130_fd_sc_hd__or2_1 _7529_ (.A(_2553_),
    .B(_2659_),
    .X(_2660_));
 sky130_fd_sc_hd__nand2_1 _7530_ (.A(net8),
    .B(net43),
    .Y(_2661_));
 sky130_fd_sc_hd__a21bo_1 _7531_ (.A1(_2553_),
    .A2(_2659_),
    .B1_N(_2661_),
    .X(_2663_));
 sky130_fd_sc_hd__nand2_1 _7532_ (.A(_2660_),
    .B(_2663_),
    .Y(_2664_));
 sky130_fd_sc_hd__a31o_1 _7533_ (.A1(_2549_),
    .A2(_2660_),
    .A3(_2663_),
    .B1(_2550_),
    .X(_2665_));
 sky130_fd_sc_hd__nor2_1 _7534_ (.A(_2544_),
    .B(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__nand2_1 _7535_ (.A(net10),
    .B(net43),
    .Y(_2667_));
 sky130_fd_sc_hd__a21boi_2 _7536_ (.A1(_2544_),
    .A2(_2665_),
    .B1_N(_2667_),
    .Y(_2668_));
 sky130_fd_sc_hd__o31ai_4 _7537_ (.A1(_2539_),
    .A2(_2666_),
    .A3(_2668_),
    .B1(_2542_),
    .Y(_2669_));
 sky130_fd_sc_hd__xnor2_1 _7538_ (.A(_2517_),
    .B(_2520_),
    .Y(_2670_));
 sky130_fd_sc_hd__xnor2_2 _7539_ (.A(_2522_),
    .B(_2670_),
    .Y(_2671_));
 sky130_fd_sc_hd__or2_1 _7540_ (.A(_2669_),
    .B(_2671_),
    .X(_2672_));
 sky130_fd_sc_hd__and2_1 _7541_ (.A(_2669_),
    .B(_2671_),
    .X(_2674_));
 sky130_fd_sc_hd__nand2_1 _7542_ (.A(net13),
    .B(net43),
    .Y(_2675_));
 sky130_fd_sc_hd__a21bo_1 _7543_ (.A1(_2669_),
    .A2(_2671_),
    .B1_N(_2675_),
    .X(_2676_));
 sky130_fd_sc_hd__o211a_1 _7544_ (.A1(_2669_),
    .A2(_2671_),
    .B1(net13),
    .C1(net43),
    .X(_2677_));
 sky130_fd_sc_hd__o31a_1 _7545_ (.A1(_2534_),
    .A2(_2674_),
    .A3(_2677_),
    .B1(_2533_),
    .X(_2678_));
 sky130_fd_sc_hd__xor2_1 _7546_ (.A(_2524_),
    .B(_2525_),
    .X(_2679_));
 sky130_fd_sc_hd__xnor2_1 _7547_ (.A(_3976_),
    .B(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__nor2_1 _7548_ (.A(_2678_),
    .B(_2680_),
    .Y(_2681_));
 sky130_fd_sc_hd__nand2_1 _7549_ (.A(net15),
    .B(net43),
    .Y(_2682_));
 sky130_fd_sc_hd__a21boi_1 _7550_ (.A1(_2678_),
    .A2(_2680_),
    .B1_N(_2682_),
    .Y(_2683_));
 sky130_fd_sc_hd__nor2_1 _7551_ (.A(_2681_),
    .B(_2683_),
    .Y(_2685_));
 sky130_fd_sc_hd__or3_1 _7552_ (.A(_2528_),
    .B(_2681_),
    .C(_2683_),
    .X(_2686_));
 sky130_fd_sc_hd__o21ai_1 _7553_ (.A1(_2681_),
    .A2(_2683_),
    .B1(_2528_),
    .Y(_2687_));
 sky130_fd_sc_hd__and3_1 _7554_ (.A(_3975_),
    .B(_2686_),
    .C(_2687_),
    .X(_2688_));
 sky130_fd_sc_hd__a21o_1 _7555_ (.A1(_2686_),
    .A2(_2687_),
    .B1(_3975_),
    .X(_2689_));
 sky130_fd_sc_hd__and2_1 _7556_ (.A(net13),
    .B(net45),
    .X(_2690_));
 sky130_fd_sc_hd__a22o_1 _7557_ (.A1(_2533_),
    .A2(_2535_),
    .B1(_2672_),
    .B2(_2676_),
    .X(_2691_));
 sky130_fd_sc_hd__nand4_1 _7558_ (.A(_2533_),
    .B(_2535_),
    .C(_2672_),
    .D(_2676_),
    .Y(_2692_));
 sky130_fd_sc_hd__a21oi_1 _7559_ (.A1(_2691_),
    .A2(_2692_),
    .B1(_2690_),
    .Y(_2693_));
 sky130_fd_sc_hd__a21o_1 _7560_ (.A1(_2691_),
    .A2(_2692_),
    .B1(_2690_),
    .X(_2694_));
 sky130_fd_sc_hd__and3_1 _7561_ (.A(_2690_),
    .B(_2691_),
    .C(_2692_),
    .X(_2696_));
 sky130_fd_sc_hd__xor2_1 _7562_ (.A(_2669_),
    .B(_2671_),
    .X(_2697_));
 sky130_fd_sc_hd__xnor2_1 _7563_ (.A(_2675_),
    .B(_2697_),
    .Y(_2698_));
 sky130_fd_sc_hd__and2_1 _7564_ (.A(net10),
    .B(net45),
    .X(_2699_));
 sky130_fd_sc_hd__o22ai_2 _7565_ (.A1(_2539_),
    .A2(_2540_),
    .B1(_2666_),
    .B2(_2668_),
    .Y(_2700_));
 sky130_fd_sc_hd__or4_1 _7566_ (.A(_2539_),
    .B(_2540_),
    .C(_2666_),
    .D(_2668_),
    .X(_2701_));
 sky130_fd_sc_hd__a21oi_1 _7567_ (.A1(_2700_),
    .A2(_2701_),
    .B1(_2699_),
    .Y(_2702_));
 sky130_fd_sc_hd__a21o_1 _7568_ (.A1(_2700_),
    .A2(_2701_),
    .B1(_2699_),
    .X(_2703_));
 sky130_fd_sc_hd__and3_1 _7569_ (.A(_2699_),
    .B(_2700_),
    .C(_2701_),
    .X(_2704_));
 sky130_fd_sc_hd__xor2_1 _7570_ (.A(_2544_),
    .B(_2665_),
    .X(_2705_));
 sky130_fd_sc_hd__xnor2_1 _7571_ (.A(_2667_),
    .B(_2705_),
    .Y(_2707_));
 sky130_fd_sc_hd__nand2_1 _7572_ (.A(net8),
    .B(net45),
    .Y(_2708_));
 sky130_fd_sc_hd__nor2_1 _7573_ (.A(_2548_),
    .B(_2550_),
    .Y(_2709_));
 sky130_fd_sc_hd__xor2_1 _7574_ (.A(_2664_),
    .B(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__nor2_1 _7575_ (.A(_2708_),
    .B(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__nand2_1 _7576_ (.A(_2708_),
    .B(_2710_),
    .Y(_2712_));
 sky130_fd_sc_hd__nand2_1 _7577_ (.A(net6),
    .B(net45),
    .Y(_2713_));
 sky130_fd_sc_hd__and2b_1 _7578_ (.A_N(_2557_),
    .B(_2558_),
    .X(_2714_));
 sky130_fd_sc_hd__xnor2_2 _7579_ (.A(_2658_),
    .B(_2714_),
    .Y(_2715_));
 sky130_fd_sc_hd__a21o_1 _7580_ (.A1(net6),
    .A2(net45),
    .B1(_2715_),
    .X(_2716_));
 sky130_fd_sc_hd__and3_1 _7581_ (.A(net6),
    .B(net45),
    .C(_2715_),
    .X(_2718_));
 sky130_fd_sc_hd__nand2_1 _7582_ (.A(net4),
    .B(net45),
    .Y(_2719_));
 sky130_fd_sc_hd__xnor2_1 _7583_ (.A(_2559_),
    .B(_2562_),
    .Y(_2720_));
 sky130_fd_sc_hd__xnor2_1 _7584_ (.A(_2649_),
    .B(_2720_),
    .Y(_2721_));
 sky130_fd_sc_hd__a21o_1 _7585_ (.A1(net4),
    .A2(net45),
    .B1(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__and3_1 _7586_ (.A(net4),
    .B(net45),
    .C(_2721_),
    .X(_2723_));
 sky130_fd_sc_hd__and2_1 _7587_ (.A(net2),
    .B(net45),
    .X(_2724_));
 sky130_fd_sc_hd__xnor2_1 _7588_ (.A(_2565_),
    .B(_2567_),
    .Y(_2725_));
 sky130_fd_sc_hd__o21bai_1 _7589_ (.A1(_2638_),
    .A2(_2642_),
    .B1_N(_2725_),
    .Y(_2726_));
 sky130_fd_sc_hd__or3b_1 _7590_ (.A(_2638_),
    .B(_2642_),
    .C_N(_2725_),
    .X(_2727_));
 sky130_fd_sc_hd__a21oi_1 _7591_ (.A1(_2726_),
    .A2(_2727_),
    .B1(_2724_),
    .Y(_2729_));
 sky130_fd_sc_hd__a21o_1 _7592_ (.A1(_2726_),
    .A2(_2727_),
    .B1(_2724_),
    .X(_2730_));
 sky130_fd_sc_hd__and3_1 _7593_ (.A(_2724_),
    .B(_2726_),
    .C(_2727_),
    .X(_2731_));
 sky130_fd_sc_hd__nand2_1 _7594_ (.A(net31),
    .B(net45),
    .Y(_2732_));
 sky130_fd_sc_hd__xor2_1 _7595_ (.A(_2570_),
    .B(_2572_),
    .X(_2733_));
 sky130_fd_sc_hd__a21o_1 _7596_ (.A1(_2631_),
    .A2(_2634_),
    .B1(_2733_),
    .X(_2734_));
 sky130_fd_sc_hd__nand3_1 _7597_ (.A(_2631_),
    .B(_2634_),
    .C(_2733_),
    .Y(_2735_));
 sky130_fd_sc_hd__a21oi_1 _7598_ (.A1(_2734_),
    .A2(_2735_),
    .B1(_2732_),
    .Y(_2736_));
 sky130_fd_sc_hd__a21o_1 _7599_ (.A1(_2734_),
    .A2(_2735_),
    .B1(_2732_),
    .X(_2737_));
 sky130_fd_sc_hd__nand3_1 _7600_ (.A(_2732_),
    .B(_2734_),
    .C(_2735_),
    .Y(_2738_));
 sky130_fd_sc_hd__and2_1 _7601_ (.A(net29),
    .B(net45),
    .X(_2740_));
 sky130_fd_sc_hd__xnor2_1 _7602_ (.A(_2576_),
    .B(_2578_),
    .Y(_2741_));
 sky130_fd_sc_hd__a21o_1 _7603_ (.A1(_2623_),
    .A2(_2625_),
    .B1(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__nand3_1 _7604_ (.A(_2623_),
    .B(_2625_),
    .C(_2741_),
    .Y(_2743_));
 sky130_fd_sc_hd__a21o_1 _7605_ (.A1(_2742_),
    .A2(_2743_),
    .B1(_2740_),
    .X(_2744_));
 sky130_fd_sc_hd__and3_1 _7606_ (.A(_2740_),
    .B(_2742_),
    .C(_2743_),
    .X(_2745_));
 sky130_fd_sc_hd__nand3_1 _7607_ (.A(_2740_),
    .B(_2742_),
    .C(_2743_),
    .Y(_2746_));
 sky130_fd_sc_hd__nand2_1 _7608_ (.A(net27),
    .B(net45),
    .Y(_2747_));
 sky130_fd_sc_hd__xor2_1 _7609_ (.A(_2581_),
    .B(_2583_),
    .X(_2748_));
 sky130_fd_sc_hd__xnor2_1 _7610_ (.A(_2619_),
    .B(_2748_),
    .Y(_2749_));
 sky130_fd_sc_hd__a21o_1 _7611_ (.A1(net27),
    .A2(net45),
    .B1(_2749_),
    .X(_2751_));
 sky130_fd_sc_hd__and3_1 _7612_ (.A(net27),
    .B(net45),
    .C(_2749_),
    .X(_2752_));
 sky130_fd_sc_hd__nand2_1 _7613_ (.A(net26),
    .B(net45),
    .Y(_2753_));
 sky130_fd_sc_hd__xor2_1 _7614_ (.A(_2587_),
    .B(_2589_),
    .X(_2754_));
 sky130_fd_sc_hd__xnor2_1 _7615_ (.A(_2617_),
    .B(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__a21o_1 _7616_ (.A1(net26),
    .A2(net45),
    .B1(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__and3_1 _7617_ (.A(net26),
    .B(net45),
    .C(_2755_),
    .X(_2757_));
 sky130_fd_sc_hd__nand2_1 _7618_ (.A(net23),
    .B(net45),
    .Y(_2758_));
 sky130_fd_sc_hd__o22ai_2 _7619_ (.A1(_2595_),
    .A2(_2597_),
    .B1(_2603_),
    .B2(_2616_),
    .Y(_2759_));
 sky130_fd_sc_hd__or4_1 _7620_ (.A(_2595_),
    .B(_2597_),
    .C(_2603_),
    .D(_2616_),
    .X(_2760_));
 sky130_fd_sc_hd__and3_1 _7621_ (.A(_2758_),
    .B(_2759_),
    .C(_2760_),
    .X(_2762_));
 sky130_fd_sc_hd__nand3_1 _7622_ (.A(_2758_),
    .B(_2759_),
    .C(_2760_),
    .Y(_2763_));
 sky130_fd_sc_hd__a21o_1 _7623_ (.A1(_2759_),
    .A2(_2760_),
    .B1(_2758_),
    .X(_2764_));
 sky130_fd_sc_hd__o211ai_1 _7624_ (.A1(_2602_),
    .A2(_2603_),
    .B1(_2608_),
    .C1(_2614_),
    .Y(_2765_));
 sky130_fd_sc_hd__a211o_1 _7625_ (.A1(_2608_),
    .A2(_2614_),
    .B1(_2602_),
    .C1(_2603_),
    .X(_2766_));
 sky130_fd_sc_hd__a22o_1 _7626_ (.A1(net12),
    .A2(net45),
    .B1(_2765_),
    .B2(_2766_),
    .X(_2767_));
 sky130_fd_sc_hd__nand4_1 _7627_ (.A(net12),
    .B(net45),
    .C(_2765_),
    .D(_2766_),
    .Y(_2768_));
 sky130_fd_sc_hd__nand2b_1 _7628_ (.A_N(_2614_),
    .B(_2608_),
    .Y(_2769_));
 sky130_fd_sc_hd__a21bo_1 _7629_ (.A1(_2608_),
    .A2(_2609_),
    .B1_N(_2613_),
    .X(_2770_));
 sky130_fd_sc_hd__and4_1 _7630_ (.A(net1),
    .B(net45),
    .C(_2769_),
    .D(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__a21boi_1 _7631_ (.A1(_2767_),
    .A2(_2771_),
    .B1_N(_2768_),
    .Y(_2773_));
 sky130_fd_sc_hd__o21ai_1 _7632_ (.A1(_2762_),
    .A2(_2773_),
    .B1(_2764_),
    .Y(_2774_));
 sky130_fd_sc_hd__a21o_1 _7633_ (.A1(_2756_),
    .A2(_2774_),
    .B1(_2757_),
    .X(_2775_));
 sky130_fd_sc_hd__a21o_1 _7634_ (.A1(_2751_),
    .A2(_2775_),
    .B1(_2752_),
    .X(_2776_));
 sky130_fd_sc_hd__xor2_1 _7635_ (.A(_2620_),
    .B(_2622_),
    .X(_2777_));
 sky130_fd_sc_hd__xnor2_1 _7636_ (.A(_2624_),
    .B(_2777_),
    .Y(_2778_));
 sky130_fd_sc_hd__or2_1 _7637_ (.A(_2776_),
    .B(_2778_),
    .X(_2779_));
 sky130_fd_sc_hd__nand2_1 _7638_ (.A(net28),
    .B(net45),
    .Y(_2780_));
 sky130_fd_sc_hd__a21bo_1 _7639_ (.A1(_2776_),
    .A2(_2778_),
    .B1_N(_2780_),
    .X(_2781_));
 sky130_fd_sc_hd__a31o_1 _7640_ (.A1(_2744_),
    .A2(_2779_),
    .A3(_2781_),
    .B1(_2745_),
    .X(_2782_));
 sky130_fd_sc_hd__xnor2_1 _7641_ (.A(_2626_),
    .B(_2628_),
    .Y(_2784_));
 sky130_fd_sc_hd__xnor2_2 _7642_ (.A(_2632_),
    .B(_2784_),
    .Y(_2785_));
 sky130_fd_sc_hd__or2_1 _7643_ (.A(_2782_),
    .B(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__and2_1 _7644_ (.A(_2782_),
    .B(_2785_),
    .X(_2787_));
 sky130_fd_sc_hd__nand2_1 _7645_ (.A(net30),
    .B(net45),
    .Y(_2788_));
 sky130_fd_sc_hd__a21bo_1 _7646_ (.A1(_2782_),
    .A2(_2785_),
    .B1_N(_2788_),
    .X(_2789_));
 sky130_fd_sc_hd__o211a_1 _7647_ (.A1(_2782_),
    .A2(_2785_),
    .B1(net30),
    .C1(net45),
    .X(_2790_));
 sky130_fd_sc_hd__o31a_1 _7648_ (.A1(_2736_),
    .A2(_2787_),
    .A3(_2790_),
    .B1(_2738_),
    .X(_2791_));
 sky130_fd_sc_hd__xnor2_1 _7649_ (.A(_2635_),
    .B(_2637_),
    .Y(_2792_));
 sky130_fd_sc_hd__xnor2_1 _7650_ (.A(_2641_),
    .B(_2792_),
    .Y(_2793_));
 sky130_fd_sc_hd__or2_1 _7651_ (.A(_2791_),
    .B(_2793_),
    .X(_2795_));
 sky130_fd_sc_hd__and2_1 _7652_ (.A(net32),
    .B(net45),
    .X(_2796_));
 sky130_fd_sc_hd__a21o_1 _7653_ (.A1(_2791_),
    .A2(_2793_),
    .B1(_2796_),
    .X(_2797_));
 sky130_fd_sc_hd__a31o_1 _7654_ (.A1(_2730_),
    .A2(_2795_),
    .A3(_2797_),
    .B1(_2731_),
    .X(_2798_));
 sky130_fd_sc_hd__and2b_1 _7655_ (.A_N(_2646_),
    .B(_2647_),
    .X(_2799_));
 sky130_fd_sc_hd__xnor2_1 _7656_ (.A(_2648_),
    .B(_2799_),
    .Y(_2800_));
 sky130_fd_sc_hd__or2_1 _7657_ (.A(_2798_),
    .B(_2800_),
    .X(_2801_));
 sky130_fd_sc_hd__nand2_1 _7658_ (.A(net3),
    .B(net45),
    .Y(_2802_));
 sky130_fd_sc_hd__a21bo_1 _7659_ (.A1(_2798_),
    .A2(_2800_),
    .B1_N(_2802_),
    .X(_2803_));
 sky130_fd_sc_hd__a31o_2 _7660_ (.A1(_2722_),
    .A2(_2801_),
    .A3(_2803_),
    .B1(_2723_),
    .X(_2804_));
 sky130_fd_sc_hd__nor2_1 _7661_ (.A(_2654_),
    .B(_2655_),
    .Y(_2806_));
 sky130_fd_sc_hd__xnor2_1 _7662_ (.A(_2656_),
    .B(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__or2_1 _7663_ (.A(_2804_),
    .B(_2807_),
    .X(_2808_));
 sky130_fd_sc_hd__nand2_1 _7664_ (.A(net5),
    .B(net45),
    .Y(_2809_));
 sky130_fd_sc_hd__a21bo_1 _7665_ (.A1(_2804_),
    .A2(_2807_),
    .B1_N(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__a31o_1 _7666_ (.A1(_2716_),
    .A2(_2808_),
    .A3(_2810_),
    .B1(_2718_),
    .X(_2811_));
 sky130_fd_sc_hd__xor2_1 _7667_ (.A(_2553_),
    .B(_2659_),
    .X(_2812_));
 sky130_fd_sc_hd__xnor2_2 _7668_ (.A(_2661_),
    .B(_2812_),
    .Y(_2813_));
 sky130_fd_sc_hd__a311o_1 _7669_ (.A1(_2716_),
    .A2(_2808_),
    .A3(_2810_),
    .B1(_2813_),
    .C1(_2718_),
    .X(_2814_));
 sky130_fd_sc_hd__and2_1 _7670_ (.A(_2811_),
    .B(_2813_),
    .X(_2815_));
 sky130_fd_sc_hd__nand2_1 _7671_ (.A(net7),
    .B(net45),
    .Y(_2817_));
 sky130_fd_sc_hd__a21bo_1 _7672_ (.A1(_2811_),
    .A2(_2813_),
    .B1_N(_2817_),
    .X(_2818_));
 sky130_fd_sc_hd__and3_1 _7673_ (.A(net7),
    .B(net45),
    .C(_2814_),
    .X(_2819_));
 sky130_fd_sc_hd__a311oi_1 _7674_ (.A1(_2712_),
    .A2(_2814_),
    .A3(_2818_),
    .B1(_2711_),
    .C1(_2707_),
    .Y(_2820_));
 sky130_fd_sc_hd__a311o_1 _7675_ (.A1(_2712_),
    .A2(_2814_),
    .A3(_2818_),
    .B1(_2711_),
    .C1(_2707_),
    .X(_2821_));
 sky130_fd_sc_hd__o311a_1 _7676_ (.A1(_2711_),
    .A2(_2815_),
    .A3(_2819_),
    .B1(_2712_),
    .C1(_2707_),
    .X(_2822_));
 sky130_fd_sc_hd__nand2_1 _7677_ (.A(net9),
    .B(net45),
    .Y(_2823_));
 sky130_fd_sc_hd__a31o_1 _7678_ (.A1(net9),
    .A2(net45),
    .A3(_2821_),
    .B1(_2822_),
    .X(_2824_));
 sky130_fd_sc_hd__a311o_1 _7679_ (.A1(net9),
    .A2(net45),
    .A3(_2821_),
    .B1(_2822_),
    .C1(_2704_),
    .X(_2825_));
 sky130_fd_sc_hd__a21o_1 _7680_ (.A1(_2703_),
    .A2(_2825_),
    .B1(_2698_),
    .X(_2826_));
 sky130_fd_sc_hd__nand3_1 _7681_ (.A(_2698_),
    .B(_2703_),
    .C(_2825_),
    .Y(_2828_));
 sky130_fd_sc_hd__and2_1 _7682_ (.A(net11),
    .B(net45),
    .X(_2829_));
 sky130_fd_sc_hd__a31o_1 _7683_ (.A1(_2698_),
    .A2(_2703_),
    .A3(_2825_),
    .B1(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__nand2_1 _7684_ (.A(_2826_),
    .B(_2830_),
    .Y(_2831_));
 sky130_fd_sc_hd__a31oi_2 _7685_ (.A1(_2694_),
    .A2(_2826_),
    .A3(_2830_),
    .B1(_2696_),
    .Y(_2832_));
 sky130_fd_sc_hd__xnor2_1 _7686_ (.A(_2678_),
    .B(_2680_),
    .Y(_2833_));
 sky130_fd_sc_hd__xnor2_1 _7687_ (.A(_2682_),
    .B(_2833_),
    .Y(_2834_));
 sky130_fd_sc_hd__and2_1 _7688_ (.A(_2832_),
    .B(_2834_),
    .X(_2835_));
 sky130_fd_sc_hd__nand2_1 _7689_ (.A(net14),
    .B(net45),
    .Y(_2836_));
 sky130_fd_sc_hd__o21a_1 _7690_ (.A1(_2832_),
    .A2(_2834_),
    .B1(_2836_),
    .X(_2837_));
 sky130_fd_sc_hd__nor2_1 _7691_ (.A(_2835_),
    .B(_2837_),
    .Y(_2839_));
 sky130_fd_sc_hd__o31ai_2 _7692_ (.A1(_2688_),
    .A2(_2835_),
    .A3(_2837_),
    .B1(_2689_),
    .Y(_2840_));
 sky130_fd_sc_hd__a22o_1 _7693_ (.A1(net43),
    .A2(_2526_),
    .B1(_2527_),
    .B2(_2685_),
    .X(_2841_));
 sky130_fd_sc_hd__o21ba_1 _7694_ (.A1(_2840_),
    .A2(_2841_),
    .B1_N(_3974_),
    .X(_2842_));
 sky130_fd_sc_hd__a21o_1 _7695_ (.A1(net46),
    .A2(_1716_),
    .B1(_2842_),
    .X(_2843_));
 sky130_fd_sc_hd__a21bo_1 _7696_ (.A1(net46),
    .A2(_2842_),
    .B1_N(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__nand2_1 _7697_ (.A(net14),
    .B(net46),
    .Y(_2845_));
 sky130_fd_sc_hd__and2b_1 _7698_ (.A_N(_2688_),
    .B(_2689_),
    .X(_2846_));
 sky130_fd_sc_hd__xor2_1 _7699_ (.A(_2839_),
    .B(_2846_),
    .X(_2847_));
 sky130_fd_sc_hd__nand2b_1 _7700_ (.A_N(_2847_),
    .B(_2845_),
    .Y(_2848_));
 sky130_fd_sc_hd__and3_1 _7701_ (.A(net14),
    .B(net46),
    .C(_2847_),
    .X(_2850_));
 sky130_fd_sc_hd__nand2_1 _7702_ (.A(net11),
    .B(net46),
    .Y(_2851_));
 sky130_fd_sc_hd__nor2_1 _7703_ (.A(_2693_),
    .B(_2696_),
    .Y(_2852_));
 sky130_fd_sc_hd__xor2_1 _7704_ (.A(_2831_),
    .B(_2852_),
    .X(_2853_));
 sky130_fd_sc_hd__and2_1 _7705_ (.A(_2851_),
    .B(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__or2_1 _7706_ (.A(_2851_),
    .B(_2853_),
    .X(_2855_));
 sky130_fd_sc_hd__nand2_1 _7707_ (.A(net9),
    .B(net46),
    .Y(_2856_));
 sky130_fd_sc_hd__nor2_1 _7708_ (.A(_2702_),
    .B(_2704_),
    .Y(_2857_));
 sky130_fd_sc_hd__xnor2_1 _7709_ (.A(_2824_),
    .B(_2857_),
    .Y(_2858_));
 sky130_fd_sc_hd__nand2_1 _7710_ (.A(_2856_),
    .B(_2858_),
    .Y(_2859_));
 sky130_fd_sc_hd__nor2_1 _7711_ (.A(_2856_),
    .B(_2858_),
    .Y(_2861_));
 sky130_fd_sc_hd__xor2_1 _7712_ (.A(_2708_),
    .B(_2710_),
    .X(_2862_));
 sky130_fd_sc_hd__or3_1 _7713_ (.A(_2815_),
    .B(_2819_),
    .C(_2862_),
    .X(_2863_));
 sky130_fd_sc_hd__o21ai_1 _7714_ (.A1(_2815_),
    .A2(_2819_),
    .B1(_2862_),
    .Y(_2864_));
 sky130_fd_sc_hd__and4_1 _7715_ (.A(net7),
    .B(net46),
    .C(_2863_),
    .D(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__a22oi_2 _7716_ (.A1(net7),
    .A2(net46),
    .B1(_2863_),
    .B2(_2864_),
    .Y(_2866_));
 sky130_fd_sc_hd__a22o_1 _7717_ (.A1(net7),
    .A2(net46),
    .B1(_2863_),
    .B2(_2864_),
    .X(_2867_));
 sky130_fd_sc_hd__nand2_1 _7718_ (.A(net5),
    .B(net46),
    .Y(_2868_));
 sky130_fd_sc_hd__xor2_1 _7719_ (.A(_2713_),
    .B(_2715_),
    .X(_2869_));
 sky130_fd_sc_hd__a21o_1 _7720_ (.A1(_2808_),
    .A2(_2810_),
    .B1(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__nand3_1 _7721_ (.A(_2808_),
    .B(_2810_),
    .C(_2869_),
    .Y(_2872_));
 sky130_fd_sc_hd__and3_1 _7722_ (.A(_2868_),
    .B(_2870_),
    .C(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__nand3_1 _7723_ (.A(_2868_),
    .B(_2870_),
    .C(_2872_),
    .Y(_2874_));
 sky130_fd_sc_hd__a21oi_1 _7724_ (.A1(_2870_),
    .A2(_2872_),
    .B1(_2868_),
    .Y(_2875_));
 sky130_fd_sc_hd__and2_1 _7725_ (.A(net3),
    .B(net46),
    .X(_2876_));
 sky130_fd_sc_hd__xnor2_1 _7726_ (.A(_2719_),
    .B(_2721_),
    .Y(_2877_));
 sky130_fd_sc_hd__a21o_1 _7727_ (.A1(_2801_),
    .A2(_2803_),
    .B1(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__nand3_1 _7728_ (.A(_2801_),
    .B(_2803_),
    .C(_2877_),
    .Y(_2879_));
 sky130_fd_sc_hd__and3_1 _7729_ (.A(_2876_),
    .B(_2878_),
    .C(_2879_),
    .X(_2880_));
 sky130_fd_sc_hd__nand3_1 _7730_ (.A(_2876_),
    .B(_2878_),
    .C(_2879_),
    .Y(_2881_));
 sky130_fd_sc_hd__a21o_1 _7731_ (.A1(_2878_),
    .A2(_2879_),
    .B1(_2876_),
    .X(_2883_));
 sky130_fd_sc_hd__and2_1 _7732_ (.A(net32),
    .B(net46),
    .X(_2884_));
 sky130_fd_sc_hd__a2bb2o_1 _7733_ (.A1_N(_2729_),
    .A2_N(_2731_),
    .B1(_2795_),
    .B2(_2797_),
    .X(_2885_));
 sky130_fd_sc_hd__or4bb_1 _7734_ (.A(_2729_),
    .B(_2731_),
    .C_N(_2795_),
    .D_N(_2797_),
    .X(_2886_));
 sky130_fd_sc_hd__a21o_1 _7735_ (.A1(_2885_),
    .A2(_2886_),
    .B1(_2884_),
    .X(_2887_));
 sky130_fd_sc_hd__and3_1 _7736_ (.A(_2884_),
    .B(_2885_),
    .C(_2886_),
    .X(_2888_));
 sky130_fd_sc_hd__nand3_1 _7737_ (.A(_2884_),
    .B(_2885_),
    .C(_2886_),
    .Y(_2889_));
 sky130_fd_sc_hd__and2_1 _7738_ (.A(net30),
    .B(net46),
    .X(_2890_));
 sky130_fd_sc_hd__a22o_1 _7739_ (.A1(_2737_),
    .A2(_2738_),
    .B1(_2786_),
    .B2(_2789_),
    .X(_2891_));
 sky130_fd_sc_hd__nand4_1 _7740_ (.A(_2737_),
    .B(_2738_),
    .C(_2786_),
    .D(_2789_),
    .Y(_2892_));
 sky130_fd_sc_hd__and3_1 _7741_ (.A(_2890_),
    .B(_2891_),
    .C(_2892_),
    .X(_2894_));
 sky130_fd_sc_hd__a21oi_1 _7742_ (.A1(_2891_),
    .A2(_2892_),
    .B1(_2890_),
    .Y(_2895_));
 sky130_fd_sc_hd__a21o_1 _7743_ (.A1(_2891_),
    .A2(_2892_),
    .B1(_2890_),
    .X(_2896_));
 sky130_fd_sc_hd__a22o_1 _7744_ (.A1(_2744_),
    .A2(_2746_),
    .B1(_2779_),
    .B2(_2781_),
    .X(_2897_));
 sky130_fd_sc_hd__nand4_1 _7745_ (.A(_2744_),
    .B(_2746_),
    .C(_2779_),
    .D(_2781_),
    .Y(_2898_));
 sky130_fd_sc_hd__and4_1 _7746_ (.A(net28),
    .B(net46),
    .C(_2897_),
    .D(_2898_),
    .X(_2899_));
 sky130_fd_sc_hd__nand4_1 _7747_ (.A(net28),
    .B(net46),
    .C(_2897_),
    .D(_2898_),
    .Y(_2900_));
 sky130_fd_sc_hd__a22o_1 _7748_ (.A1(net28),
    .A2(net46),
    .B1(_2897_),
    .B2(_2898_),
    .X(_2901_));
 sky130_fd_sc_hd__nand2_1 _7749_ (.A(net26),
    .B(net46),
    .Y(_2902_));
 sky130_fd_sc_hd__xor2_1 _7750_ (.A(_2747_),
    .B(_2749_),
    .X(_2903_));
 sky130_fd_sc_hd__xnor2_1 _7751_ (.A(_2775_),
    .B(_2903_),
    .Y(_2905_));
 sky130_fd_sc_hd__nand2b_1 _7752_ (.A_N(_2902_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__and2b_1 _7753_ (.A_N(_2905_),
    .B(_2902_),
    .X(_2907_));
 sky130_fd_sc_hd__nand2_1 _7754_ (.A(net23),
    .B(net46),
    .Y(_2908_));
 sky130_fd_sc_hd__xnor2_1 _7755_ (.A(_2753_),
    .B(_2755_),
    .Y(_2909_));
 sky130_fd_sc_hd__xnor2_1 _7756_ (.A(_2774_),
    .B(_2909_),
    .Y(_2910_));
 sky130_fd_sc_hd__nand2_1 _7757_ (.A(_2908_),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__nor2_1 _7758_ (.A(_2908_),
    .B(_2910_),
    .Y(_2912_));
 sky130_fd_sc_hd__and2_1 _7759_ (.A(net12),
    .B(net46),
    .X(_2913_));
 sky130_fd_sc_hd__and3_1 _7760_ (.A(_2763_),
    .B(_2764_),
    .C(_2773_),
    .X(_2914_));
 sky130_fd_sc_hd__a21oi_1 _7761_ (.A1(_2763_),
    .A2(_2764_),
    .B1(_2773_),
    .Y(_2916_));
 sky130_fd_sc_hd__or2_1 _7762_ (.A(_2914_),
    .B(_2916_),
    .X(_2917_));
 sky130_fd_sc_hd__and3_1 _7763_ (.A(_2767_),
    .B(_2768_),
    .C(_2771_),
    .X(_2918_));
 sky130_fd_sc_hd__a21o_1 _7764_ (.A1(_2767_),
    .A2(_2768_),
    .B1(_2771_),
    .X(_2919_));
 sky130_fd_sc_hd__and4b_1 _7765_ (.A_N(_2918_),
    .B(_2919_),
    .C(net1),
    .D(net46),
    .X(_2920_));
 sky130_fd_sc_hd__o31a_1 _7766_ (.A1(_2913_),
    .A2(_2914_),
    .A3(_2916_),
    .B1(_2920_),
    .X(_2921_));
 sky130_fd_sc_hd__a21o_1 _7767_ (.A1(_2913_),
    .A2(_2917_),
    .B1(_2921_),
    .X(_2922_));
 sky130_fd_sc_hd__a21oi_1 _7768_ (.A1(_2911_),
    .A2(_2922_),
    .B1(_2912_),
    .Y(_2923_));
 sky130_fd_sc_hd__a21oi_1 _7769_ (.A1(_2906_),
    .A2(_2923_),
    .B1(_2907_),
    .Y(_2924_));
 sky130_fd_sc_hd__xor2_1 _7770_ (.A(_2776_),
    .B(_2778_),
    .X(_2925_));
 sky130_fd_sc_hd__xnor2_1 _7771_ (.A(_2780_),
    .B(_2925_),
    .Y(_2927_));
 sky130_fd_sc_hd__or2_1 _7772_ (.A(_2924_),
    .B(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__nand2_1 _7773_ (.A(net27),
    .B(net46),
    .Y(_2929_));
 sky130_fd_sc_hd__a21bo_1 _7774_ (.A1(_2924_),
    .A2(_2927_),
    .B1_N(_2929_),
    .X(_2930_));
 sky130_fd_sc_hd__a31o_1 _7775_ (.A1(_2901_),
    .A2(_2928_),
    .A3(_2930_),
    .B1(_2899_),
    .X(_2931_));
 sky130_fd_sc_hd__xor2_1 _7776_ (.A(_2782_),
    .B(_2785_),
    .X(_2932_));
 sky130_fd_sc_hd__xnor2_2 _7777_ (.A(_2788_),
    .B(_2932_),
    .Y(_2933_));
 sky130_fd_sc_hd__or2_1 _7778_ (.A(_2931_),
    .B(_2933_),
    .X(_2934_));
 sky130_fd_sc_hd__and2_1 _7779_ (.A(_2931_),
    .B(_2933_),
    .X(_2935_));
 sky130_fd_sc_hd__and2_1 _7780_ (.A(net29),
    .B(net46),
    .X(_2936_));
 sky130_fd_sc_hd__a21o_1 _7781_ (.A1(_2931_),
    .A2(_2933_),
    .B1(_2936_),
    .X(_2938_));
 sky130_fd_sc_hd__o211a_1 _7782_ (.A1(_2931_),
    .A2(_2933_),
    .B1(net29),
    .C1(net46),
    .X(_2939_));
 sky130_fd_sc_hd__o31a_1 _7783_ (.A1(_2894_),
    .A2(_2935_),
    .A3(_2939_),
    .B1(_2896_),
    .X(_2940_));
 sky130_fd_sc_hd__xnor2_1 _7784_ (.A(_2791_),
    .B(_2793_),
    .Y(_2941_));
 sky130_fd_sc_hd__xnor2_1 _7785_ (.A(_2796_),
    .B(_2941_),
    .Y(_2942_));
 sky130_fd_sc_hd__or2_1 _7786_ (.A(_2940_),
    .B(_2942_),
    .X(_2943_));
 sky130_fd_sc_hd__and2_1 _7787_ (.A(net31),
    .B(net46),
    .X(_2944_));
 sky130_fd_sc_hd__a21o_1 _7788_ (.A1(_2940_),
    .A2(_2942_),
    .B1(_2944_),
    .X(_2945_));
 sky130_fd_sc_hd__a31o_1 _7789_ (.A1(_2887_),
    .A2(_2943_),
    .A3(_2945_),
    .B1(_2888_),
    .X(_2946_));
 sky130_fd_sc_hd__xor2_1 _7790_ (.A(_2798_),
    .B(_2800_),
    .X(_2947_));
 sky130_fd_sc_hd__xnor2_2 _7791_ (.A(_2802_),
    .B(_2947_),
    .Y(_2949_));
 sky130_fd_sc_hd__nor2_1 _7792_ (.A(_2946_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__and2_1 _7793_ (.A(_2946_),
    .B(_2949_),
    .X(_2951_));
 sky130_fd_sc_hd__and2_1 _7794_ (.A(net2),
    .B(net46),
    .X(_2952_));
 sky130_fd_sc_hd__a21oi_1 _7795_ (.A1(_2946_),
    .A2(_2949_),
    .B1(_2952_),
    .Y(_2953_));
 sky130_fd_sc_hd__o211a_1 _7796_ (.A1(_2946_),
    .A2(_2949_),
    .B1(net2),
    .C1(net46),
    .X(_2954_));
 sky130_fd_sc_hd__o31a_2 _7797_ (.A1(_2880_),
    .A2(_2951_),
    .A3(_2954_),
    .B1(_2883_),
    .X(_2955_));
 sky130_fd_sc_hd__xor2_1 _7798_ (.A(_2804_),
    .B(_2807_),
    .X(_2956_));
 sky130_fd_sc_hd__xnor2_1 _7799_ (.A(_2809_),
    .B(_2956_),
    .Y(_2957_));
 sky130_fd_sc_hd__or2_1 _7800_ (.A(_2955_),
    .B(_2957_),
    .X(_2958_));
 sky130_fd_sc_hd__and2_1 _7801_ (.A(net4),
    .B(net46),
    .X(_2960_));
 sky130_fd_sc_hd__a21o_1 _7802_ (.A1(_2955_),
    .A2(_2957_),
    .B1(_2960_),
    .X(_2961_));
 sky130_fd_sc_hd__a31o_1 _7803_ (.A1(_2874_),
    .A2(_2958_),
    .A3(_2961_),
    .B1(_2875_),
    .X(_2962_));
 sky130_fd_sc_hd__xor2_1 _7804_ (.A(_2811_),
    .B(_2813_),
    .X(_2963_));
 sky130_fd_sc_hd__xnor2_1 _7805_ (.A(_2817_),
    .B(_2963_),
    .Y(_2964_));
 sky130_fd_sc_hd__or2_1 _7806_ (.A(_2962_),
    .B(_2964_),
    .X(_2965_));
 sky130_fd_sc_hd__nand2_1 _7807_ (.A(net6),
    .B(net46),
    .Y(_2966_));
 sky130_fd_sc_hd__a21bo_1 _7808_ (.A1(_2962_),
    .A2(_2964_),
    .B1_N(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__a31o_1 _7809_ (.A1(_2867_),
    .A2(_2965_),
    .A3(_2967_),
    .B1(_2865_),
    .X(_2968_));
 sky130_fd_sc_hd__nor2_1 _7810_ (.A(_2820_),
    .B(_2822_),
    .Y(_2969_));
 sky130_fd_sc_hd__xnor2_1 _7811_ (.A(_2823_),
    .B(_2969_),
    .Y(_2971_));
 sky130_fd_sc_hd__or2_1 _7812_ (.A(_2968_),
    .B(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__and2_1 _7813_ (.A(net8),
    .B(net46),
    .X(_2973_));
 sky130_fd_sc_hd__a21o_1 _7814_ (.A1(_2968_),
    .A2(_2971_),
    .B1(_2973_),
    .X(_2974_));
 sky130_fd_sc_hd__a31o_1 _7815_ (.A1(_2859_),
    .A2(_2972_),
    .A3(_2974_),
    .B1(_2861_),
    .X(_2975_));
 sky130_fd_sc_hd__and2_1 _7816_ (.A(_2826_),
    .B(_2828_),
    .X(_2976_));
 sky130_fd_sc_hd__xor2_2 _7817_ (.A(_2829_),
    .B(_2976_),
    .X(_2977_));
 sky130_fd_sc_hd__nor2_1 _7818_ (.A(_2975_),
    .B(_2977_),
    .Y(_2978_));
 sky130_fd_sc_hd__nand2_1 _7819_ (.A(_2975_),
    .B(_2977_),
    .Y(_2979_));
 sky130_fd_sc_hd__and2_1 _7820_ (.A(net10),
    .B(net46),
    .X(_2980_));
 sky130_fd_sc_hd__a21oi_1 _7821_ (.A1(_2975_),
    .A2(_2977_),
    .B1(_2980_),
    .Y(_2982_));
 sky130_fd_sc_hd__o211ai_1 _7822_ (.A1(_2975_),
    .A2(_2977_),
    .B1(net10),
    .C1(net46),
    .Y(_2983_));
 sky130_fd_sc_hd__xnor2_1 _7823_ (.A(_2832_),
    .B(_2834_),
    .Y(_2984_));
 sky130_fd_sc_hd__xnor2_1 _7824_ (.A(_2836_),
    .B(_2984_),
    .Y(_2985_));
 sky130_fd_sc_hd__o311a_1 _7825_ (.A1(_2854_),
    .A2(_2978_),
    .A3(_2982_),
    .B1(_2985_),
    .C1(_2855_),
    .X(_2986_));
 sky130_fd_sc_hd__a311o_1 _7826_ (.A1(_2855_),
    .A2(_2979_),
    .A3(_2983_),
    .B1(_2985_),
    .C1(_2854_),
    .X(_2987_));
 sky130_fd_sc_hd__inv_2 _7827_ (.A(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__nand2_1 _7828_ (.A(net13),
    .B(net46),
    .Y(_2989_));
 sky130_fd_sc_hd__and3b_1 _7829_ (.A_N(_2986_),
    .B(net46),
    .C(net13),
    .X(_2990_));
 sky130_fd_sc_hd__a21oi_1 _7830_ (.A1(_2987_),
    .A2(_2989_),
    .B1(_2986_),
    .Y(_2991_));
 sky130_fd_sc_hd__xnor2_1 _7831_ (.A(_2840_),
    .B(_2841_),
    .Y(_2993_));
 sky130_fd_sc_hd__xor2_1 _7832_ (.A(_3974_),
    .B(_2993_),
    .X(_2994_));
 sky130_fd_sc_hd__a211oi_1 _7833_ (.A1(_2848_),
    .A2(_2991_),
    .B1(_2994_),
    .C1(_2850_),
    .Y(_2995_));
 sky130_fd_sc_hd__o311a_1 _7834_ (.A1(_2850_),
    .A2(_2988_),
    .A3(_2990_),
    .B1(_2994_),
    .C1(_2848_),
    .X(_2996_));
 sky130_fd_sc_hd__nand2_1 _7835_ (.A(net15),
    .B(net46),
    .Y(_2997_));
 sky130_fd_sc_hd__o21bai_1 _7836_ (.A1(_2995_),
    .A2(_2997_),
    .B1_N(_2996_),
    .Y(_2998_));
 sky130_fd_sc_hd__xnor2_1 _7837_ (.A(_2844_),
    .B(_2998_),
    .Y(_2999_));
 sky130_fd_sc_hd__a21oi_1 _7838_ (.A1(net15),
    .A2(net47),
    .B1(_2999_),
    .Y(_3000_));
 sky130_fd_sc_hd__nand3_1 _7839_ (.A(net15),
    .B(net47),
    .C(_2999_),
    .Y(_3001_));
 sky130_fd_sc_hd__xor2_1 _7840_ (.A(_2845_),
    .B(_2847_),
    .X(_3002_));
 sky130_fd_sc_hd__xnor2_1 _7841_ (.A(_2991_),
    .B(_3002_),
    .Y(_3004_));
 sky130_fd_sc_hd__a21oi_1 _7842_ (.A1(net13),
    .A2(net47),
    .B1(_3004_),
    .Y(_3005_));
 sky130_fd_sc_hd__or3b_1 _7843_ (.A(_0000_),
    .B(_0110_),
    .C_N(_3004_),
    .X(_3006_));
 sky130_fd_sc_hd__and2_1 _7844_ (.A(net10),
    .B(net47),
    .X(_3007_));
 sky130_fd_sc_hd__xor2_1 _7845_ (.A(_2851_),
    .B(_2853_),
    .X(_3008_));
 sky130_fd_sc_hd__o21bai_1 _7846_ (.A1(_2978_),
    .A2(_2982_),
    .B1_N(_3008_),
    .Y(_3009_));
 sky130_fd_sc_hd__or3b_1 _7847_ (.A(_2978_),
    .B(_2982_),
    .C_N(_3008_),
    .X(_3010_));
 sky130_fd_sc_hd__a21oi_1 _7848_ (.A1(_3009_),
    .A2(_3010_),
    .B1(_3007_),
    .Y(_3011_));
 sky130_fd_sc_hd__a21o_1 _7849_ (.A1(_3009_),
    .A2(_3010_),
    .B1(_3007_),
    .X(_3012_));
 sky130_fd_sc_hd__and3_1 _7850_ (.A(_3007_),
    .B(_3009_),
    .C(_3010_),
    .X(_3013_));
 sky130_fd_sc_hd__and2_1 _7851_ (.A(net8),
    .B(net47),
    .X(_3015_));
 sky130_fd_sc_hd__xor2_1 _7852_ (.A(_2856_),
    .B(_2858_),
    .X(_3016_));
 sky130_fd_sc_hd__a21o_1 _7853_ (.A1(_2972_),
    .A2(_2974_),
    .B1(_3016_),
    .X(_3017_));
 sky130_fd_sc_hd__nand3_1 _7854_ (.A(_2972_),
    .B(_2974_),
    .C(_3016_),
    .Y(_3018_));
 sky130_fd_sc_hd__a21oi_1 _7855_ (.A1(_3017_),
    .A2(_3018_),
    .B1(_3015_),
    .Y(_3019_));
 sky130_fd_sc_hd__a21o_1 _7856_ (.A1(_3017_),
    .A2(_3018_),
    .B1(_3015_),
    .X(_3020_));
 sky130_fd_sc_hd__and3_1 _7857_ (.A(_3015_),
    .B(_3017_),
    .C(_3018_),
    .X(_3021_));
 sky130_fd_sc_hd__nand2_1 _7858_ (.A(net6),
    .B(net47),
    .Y(_3022_));
 sky130_fd_sc_hd__o211ai_2 _7859_ (.A1(_2865_),
    .A2(_2866_),
    .B1(_2965_),
    .C1(_2967_),
    .Y(_3023_));
 sky130_fd_sc_hd__a211o_1 _7860_ (.A1(_2965_),
    .A2(_2967_),
    .B1(_2865_),
    .C1(_2866_),
    .X(_3024_));
 sky130_fd_sc_hd__a21oi_1 _7861_ (.A1(_3023_),
    .A2(_3024_),
    .B1(_3022_),
    .Y(_3026_));
 sky130_fd_sc_hd__a21o_1 _7862_ (.A1(_3023_),
    .A2(_3024_),
    .B1(_3022_),
    .X(_3027_));
 sky130_fd_sc_hd__and3_1 _7863_ (.A(_3022_),
    .B(_3023_),
    .C(_3024_),
    .X(_3028_));
 sky130_fd_sc_hd__and2_1 _7864_ (.A(net4),
    .B(net47),
    .X(_3029_));
 sky130_fd_sc_hd__a2bb2o_1 _7865_ (.A1_N(_2873_),
    .A2_N(_2875_),
    .B1(_2958_),
    .B2(_2961_),
    .X(_3030_));
 sky130_fd_sc_hd__or4bb_1 _7866_ (.A(_2873_),
    .B(_2875_),
    .C_N(_2958_),
    .D_N(_2961_),
    .X(_3031_));
 sky130_fd_sc_hd__and2_1 _7867_ (.A(_3030_),
    .B(_3031_),
    .X(_3032_));
 sky130_fd_sc_hd__nor2_1 _7868_ (.A(_3029_),
    .B(_3032_),
    .Y(_3033_));
 sky130_fd_sc_hd__a21o_1 _7869_ (.A1(_3030_),
    .A2(_3031_),
    .B1(_3029_),
    .X(_3034_));
 sky130_fd_sc_hd__and3_1 _7870_ (.A(_3029_),
    .B(_3030_),
    .C(_3031_),
    .X(_3035_));
 sky130_fd_sc_hd__nand2_1 _7871_ (.A(net2),
    .B(net47),
    .Y(_3037_));
 sky130_fd_sc_hd__a211o_1 _7872_ (.A1(_2881_),
    .A2(_2883_),
    .B1(_2950_),
    .C1(_2953_),
    .X(_3038_));
 sky130_fd_sc_hd__o211ai_1 _7873_ (.A1(_2950_),
    .A2(_2953_),
    .B1(_2881_),
    .C1(_2883_),
    .Y(_3039_));
 sky130_fd_sc_hd__and3_1 _7874_ (.A(_3037_),
    .B(_3038_),
    .C(_3039_),
    .X(_3040_));
 sky130_fd_sc_hd__a21o_1 _7875_ (.A1(_3038_),
    .A2(_3039_),
    .B1(_3037_),
    .X(_3041_));
 sky130_fd_sc_hd__and2_1 _7876_ (.A(net31),
    .B(net47),
    .X(_3042_));
 sky130_fd_sc_hd__a22o_1 _7877_ (.A1(_2887_),
    .A2(_2889_),
    .B1(_2943_),
    .B2(_2945_),
    .X(_3043_));
 sky130_fd_sc_hd__nand4_1 _7878_ (.A(_2887_),
    .B(_2889_),
    .C(_2943_),
    .D(_2945_),
    .Y(_3044_));
 sky130_fd_sc_hd__and3_1 _7879_ (.A(_3042_),
    .B(_3043_),
    .C(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__a21o_1 _7880_ (.A1(_3043_),
    .A2(_3044_),
    .B1(_3042_),
    .X(_3046_));
 sky130_fd_sc_hd__and2_1 _7881_ (.A(net29),
    .B(net47),
    .X(_3048_));
 sky130_fd_sc_hd__a211oi_1 _7882_ (.A1(_2934_),
    .A2(_2938_),
    .B1(_2894_),
    .C1(_2895_),
    .Y(_3049_));
 sky130_fd_sc_hd__o211a_1 _7883_ (.A1(_2894_),
    .A2(_2895_),
    .B1(_2934_),
    .C1(_2938_),
    .X(_3050_));
 sky130_fd_sc_hd__or2_1 _7884_ (.A(_3049_),
    .B(_3050_),
    .X(_3051_));
 sky130_fd_sc_hd__or3_1 _7885_ (.A(_3048_),
    .B(_3049_),
    .C(_3050_),
    .X(_3052_));
 sky130_fd_sc_hd__o21a_1 _7886_ (.A1(_3049_),
    .A2(_3050_),
    .B1(_3048_),
    .X(_3053_));
 sky130_fd_sc_hd__nor2_1 _7887_ (.A(_4187_),
    .B(_0110_),
    .Y(_3054_));
 sky130_fd_sc_hd__a22o_1 _7888_ (.A1(_2900_),
    .A2(_2901_),
    .B1(_2928_),
    .B2(_2930_),
    .X(_3055_));
 sky130_fd_sc_hd__nand4_1 _7889_ (.A(_2900_),
    .B(_2901_),
    .C(_2928_),
    .D(_2930_),
    .Y(_3056_));
 sky130_fd_sc_hd__a21oi_1 _7890_ (.A1(_3055_),
    .A2(_3056_),
    .B1(_3054_),
    .Y(_3057_));
 sky130_fd_sc_hd__a21o_1 _7891_ (.A1(_3055_),
    .A2(_3056_),
    .B1(_3054_),
    .X(_3059_));
 sky130_fd_sc_hd__and3_1 _7892_ (.A(_3054_),
    .B(_3055_),
    .C(_3056_),
    .X(_3060_));
 sky130_fd_sc_hd__nand2_1 _7893_ (.A(net23),
    .B(net47),
    .Y(_3061_));
 sky130_fd_sc_hd__xnor2_1 _7894_ (.A(_2902_),
    .B(_2905_),
    .Y(_3062_));
 sky130_fd_sc_hd__xnor2_1 _7895_ (.A(_2923_),
    .B(_3062_),
    .Y(_3063_));
 sky130_fd_sc_hd__nand2b_1 _7896_ (.A_N(_3061_),
    .B(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__a21oi_1 _7897_ (.A1(net23),
    .A2(net47),
    .B1(_3063_),
    .Y(_3065_));
 sky130_fd_sc_hd__and2_1 _7898_ (.A(net12),
    .B(net47),
    .X(_3066_));
 sky130_fd_sc_hd__xnor2_1 _7899_ (.A(_2908_),
    .B(_2910_),
    .Y(_3067_));
 sky130_fd_sc_hd__xnor2_1 _7900_ (.A(_2922_),
    .B(_3067_),
    .Y(_3068_));
 sky130_fd_sc_hd__nor2_1 _7901_ (.A(_3066_),
    .B(_3068_),
    .Y(_3070_));
 sky130_fd_sc_hd__or2_1 _7902_ (.A(_3066_),
    .B(_3068_),
    .X(_3071_));
 sky130_fd_sc_hd__and2_1 _7903_ (.A(_3066_),
    .B(_3068_),
    .X(_3072_));
 sky130_fd_sc_hd__xor2_1 _7904_ (.A(_2913_),
    .B(_2917_),
    .X(_3073_));
 sky130_fd_sc_hd__o211ai_1 _7905_ (.A1(_2920_),
    .A2(_3073_),
    .B1(net1),
    .C1(net47),
    .Y(_3074_));
 sky130_fd_sc_hd__a21oi_1 _7906_ (.A1(_2920_),
    .A2(_3073_),
    .B1(_3074_),
    .Y(_3075_));
 sky130_fd_sc_hd__a21oi_1 _7907_ (.A1(_3071_),
    .A2(_3075_),
    .B1(_3072_),
    .Y(_3076_));
 sky130_fd_sc_hd__a21oi_1 _7908_ (.A1(_3064_),
    .A2(_3076_),
    .B1(_3065_),
    .Y(_3077_));
 sky130_fd_sc_hd__xor2_1 _7909_ (.A(_2924_),
    .B(_2927_),
    .X(_3078_));
 sky130_fd_sc_hd__xnor2_1 _7910_ (.A(_2929_),
    .B(_3078_),
    .Y(_3079_));
 sky130_fd_sc_hd__or2_1 _7911_ (.A(_3077_),
    .B(_3079_),
    .X(_3081_));
 sky130_fd_sc_hd__nand2_1 _7912_ (.A(net26),
    .B(net47),
    .Y(_3082_));
 sky130_fd_sc_hd__a21bo_1 _7913_ (.A1(_3077_),
    .A2(_3079_),
    .B1_N(_3082_),
    .X(_3083_));
 sky130_fd_sc_hd__nand2_1 _7914_ (.A(_3081_),
    .B(_3083_),
    .Y(_3084_));
 sky130_fd_sc_hd__a31o_1 _7915_ (.A1(_3059_),
    .A2(_3081_),
    .A3(_3083_),
    .B1(_3060_),
    .X(_3085_));
 sky130_fd_sc_hd__xnor2_1 _7916_ (.A(_2931_),
    .B(_2933_),
    .Y(_3086_));
 sky130_fd_sc_hd__xnor2_1 _7917_ (.A(_2936_),
    .B(_3086_),
    .Y(_3087_));
 sky130_fd_sc_hd__and2_1 _7918_ (.A(_3085_),
    .B(_3087_),
    .X(_3088_));
 sky130_fd_sc_hd__nand2_1 _7919_ (.A(net28),
    .B(net47),
    .Y(_3089_));
 sky130_fd_sc_hd__o211a_1 _7920_ (.A1(_3085_),
    .A2(_3087_),
    .B1(net28),
    .C1(net47),
    .X(_3090_));
 sky130_fd_sc_hd__nor2_1 _7921_ (.A(_3088_),
    .B(_3090_),
    .Y(_3092_));
 sky130_fd_sc_hd__o31a_1 _7922_ (.A1(_3053_),
    .A2(_3088_),
    .A3(_3090_),
    .B1(_3052_),
    .X(_3093_));
 sky130_fd_sc_hd__xnor2_1 _7923_ (.A(_2940_),
    .B(_2942_),
    .Y(_3094_));
 sky130_fd_sc_hd__xnor2_1 _7924_ (.A(_2944_),
    .B(_3094_),
    .Y(_3095_));
 sky130_fd_sc_hd__or2_1 _7925_ (.A(_3093_),
    .B(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__and2_1 _7926_ (.A(net30),
    .B(net47),
    .X(_3097_));
 sky130_fd_sc_hd__a21o_1 _7927_ (.A1(_3093_),
    .A2(_3095_),
    .B1(_3097_),
    .X(_3098_));
 sky130_fd_sc_hd__nand2_1 _7928_ (.A(_3096_),
    .B(_3098_),
    .Y(_3099_));
 sky130_fd_sc_hd__a31o_1 _7929_ (.A1(_3046_),
    .A2(_3096_),
    .A3(_3098_),
    .B1(_3045_),
    .X(_3100_));
 sky130_fd_sc_hd__xnor2_1 _7930_ (.A(_2946_),
    .B(_2949_),
    .Y(_3101_));
 sky130_fd_sc_hd__xnor2_2 _7931_ (.A(_2952_),
    .B(_3101_),
    .Y(_3103_));
 sky130_fd_sc_hd__nand2_1 _7932_ (.A(_3100_),
    .B(_3103_),
    .Y(_3104_));
 sky130_fd_sc_hd__nand2_1 _7933_ (.A(net32),
    .B(net47),
    .Y(_3105_));
 sky130_fd_sc_hd__o211ai_2 _7934_ (.A1(_3100_),
    .A2(_3103_),
    .B1(net32),
    .C1(net47),
    .Y(_3106_));
 sky130_fd_sc_hd__nand2_1 _7935_ (.A(_3104_),
    .B(_3106_),
    .Y(_3107_));
 sky130_fd_sc_hd__a31oi_4 _7936_ (.A1(_3041_),
    .A2(_3104_),
    .A3(_3106_),
    .B1(_3040_),
    .Y(_3108_));
 sky130_fd_sc_hd__xnor2_1 _7937_ (.A(_2955_),
    .B(_2957_),
    .Y(_3109_));
 sky130_fd_sc_hd__xnor2_1 _7938_ (.A(_2960_),
    .B(_3109_),
    .Y(_3110_));
 sky130_fd_sc_hd__or2_1 _7939_ (.A(_3108_),
    .B(_3110_),
    .X(_3111_));
 sky130_fd_sc_hd__nand2_1 _7940_ (.A(net3),
    .B(net47),
    .Y(_3112_));
 sky130_fd_sc_hd__a21bo_1 _7941_ (.A1(_3108_),
    .A2(_3110_),
    .B1_N(_3112_),
    .X(_3114_));
 sky130_fd_sc_hd__nand2_1 _7942_ (.A(_3111_),
    .B(_3114_),
    .Y(_3115_));
 sky130_fd_sc_hd__a21oi_1 _7943_ (.A1(_3111_),
    .A2(_3114_),
    .B1(_3035_),
    .Y(_3116_));
 sky130_fd_sc_hd__a31o_1 _7944_ (.A1(_3034_),
    .A2(_3111_),
    .A3(_3114_),
    .B1(_3035_),
    .X(_3117_));
 sky130_fd_sc_hd__xnor2_1 _7945_ (.A(_2962_),
    .B(_2964_),
    .Y(_3118_));
 sky130_fd_sc_hd__xnor2_1 _7946_ (.A(_2966_),
    .B(_3118_),
    .Y(_3119_));
 sky130_fd_sc_hd__and2b_1 _7947_ (.A_N(_3117_),
    .B(_3119_),
    .X(_3120_));
 sky130_fd_sc_hd__nand2_1 _7948_ (.A(net5),
    .B(net47),
    .Y(_3121_));
 sky130_fd_sc_hd__o31a_1 _7949_ (.A1(_3033_),
    .A2(_3116_),
    .A3(_3119_),
    .B1(_3121_),
    .X(_3122_));
 sky130_fd_sc_hd__or2_1 _7950_ (.A(_3120_),
    .B(_3122_),
    .X(_3123_));
 sky130_fd_sc_hd__o31ai_2 _7951_ (.A1(_3028_),
    .A2(_3120_),
    .A3(_3122_),
    .B1(_3027_),
    .Y(_3125_));
 sky130_fd_sc_hd__xnor2_1 _7952_ (.A(_2968_),
    .B(_2971_),
    .Y(_3126_));
 sky130_fd_sc_hd__xnor2_1 _7953_ (.A(_2973_),
    .B(_3126_),
    .Y(_3127_));
 sky130_fd_sc_hd__or2_1 _7954_ (.A(_3125_),
    .B(_3127_),
    .X(_3128_));
 sky130_fd_sc_hd__nand2_1 _7955_ (.A(net7),
    .B(net47),
    .Y(_3129_));
 sky130_fd_sc_hd__a21bo_1 _7956_ (.A1(_3125_),
    .A2(_3127_),
    .B1_N(_3129_),
    .X(_3130_));
 sky130_fd_sc_hd__nand2_1 _7957_ (.A(_3128_),
    .B(_3130_),
    .Y(_3131_));
 sky130_fd_sc_hd__a21oi_1 _7958_ (.A1(_3128_),
    .A2(_3130_),
    .B1(_3021_),
    .Y(_3132_));
 sky130_fd_sc_hd__a31o_1 _7959_ (.A1(_3020_),
    .A2(_3128_),
    .A3(_3130_),
    .B1(_3021_),
    .X(_3133_));
 sky130_fd_sc_hd__xor2_1 _7960_ (.A(_2975_),
    .B(_2977_),
    .X(_3134_));
 sky130_fd_sc_hd__xnor2_1 _7961_ (.A(_2980_),
    .B(_3134_),
    .Y(_3136_));
 sky130_fd_sc_hd__nand2b_1 _7962_ (.A_N(_3133_),
    .B(_3136_),
    .Y(_3137_));
 sky130_fd_sc_hd__nand2_1 _7963_ (.A(net9),
    .B(net47),
    .Y(_3138_));
 sky130_fd_sc_hd__o31ai_1 _7964_ (.A1(_3019_),
    .A2(_3132_),
    .A3(_3136_),
    .B1(_3138_),
    .Y(_3139_));
 sky130_fd_sc_hd__nand2_1 _7965_ (.A(_3137_),
    .B(_3139_),
    .Y(_3140_));
 sky130_fd_sc_hd__a31o_1 _7966_ (.A1(_3012_),
    .A2(_3137_),
    .A3(_3139_),
    .B1(_3013_),
    .X(_3141_));
 sky130_fd_sc_hd__and2b_1 _7967_ (.A_N(_2986_),
    .B(_2987_),
    .X(_3142_));
 sky130_fd_sc_hd__xnor2_1 _7968_ (.A(_2989_),
    .B(_3142_),
    .Y(_3143_));
 sky130_fd_sc_hd__nor2_1 _7969_ (.A(_3141_),
    .B(_3143_),
    .Y(_3144_));
 sky130_fd_sc_hd__nand2_1 _7970_ (.A(net11),
    .B(net47),
    .Y(_3145_));
 sky130_fd_sc_hd__a21boi_1 _7971_ (.A1(_3141_),
    .A2(_3143_),
    .B1_N(_3145_),
    .Y(_3147_));
 sky130_fd_sc_hd__nor2_1 _7972_ (.A(_3144_),
    .B(_3147_),
    .Y(_3148_));
 sky130_fd_sc_hd__o31ai_2 _7973_ (.A1(_3005_),
    .A2(_3144_),
    .A3(_3147_),
    .B1(_3006_),
    .Y(_3149_));
 sky130_fd_sc_hd__nor2_1 _7974_ (.A(_2995_),
    .B(_2996_),
    .Y(_3150_));
 sky130_fd_sc_hd__xnor2_1 _7975_ (.A(_2997_),
    .B(_3150_),
    .Y(_3151_));
 sky130_fd_sc_hd__nor2_1 _7976_ (.A(_3149_),
    .B(_3151_),
    .Y(_3152_));
 sky130_fd_sc_hd__nand2_1 _7977_ (.A(net14),
    .B(net47),
    .Y(_3153_));
 sky130_fd_sc_hd__a21boi_1 _7978_ (.A1(_3149_),
    .A2(_3151_),
    .B1_N(_3153_),
    .Y(_3154_));
 sky130_fd_sc_hd__nor2_1 _7979_ (.A(_3152_),
    .B(_3154_),
    .Y(_3155_));
 sky130_fd_sc_hd__o31a_1 _7980_ (.A1(_3000_),
    .A2(_3152_),
    .A3(_3154_),
    .B1(_3001_),
    .X(_3156_));
 sky130_fd_sc_hd__a22oi_2 _7981_ (.A1(net46),
    .A2(_2842_),
    .B1(_2843_),
    .B2(_2998_),
    .Y(_3158_));
 sky130_fd_sc_hd__a21oi_2 _7982_ (.A1(_3156_),
    .A2(_3158_),
    .B1(_3973_),
    .Y(_3159_));
 sky130_fd_sc_hd__a21o_1 _7983_ (.A1(_1716_),
    .A2(_1760_),
    .B1(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__nand2_1 _7984_ (.A(_1760_),
    .B(_3159_),
    .Y(_3161_));
 sky130_fd_sc_hd__and2_1 _7985_ (.A(net15),
    .B(_1760_),
    .X(_3162_));
 sky130_fd_sc_hd__xor2_1 _7986_ (.A(_3156_),
    .B(_3158_),
    .X(_3163_));
 sky130_fd_sc_hd__xnor2_1 _7987_ (.A(_3973_),
    .B(_3163_),
    .Y(_3164_));
 sky130_fd_sc_hd__or2_1 _7988_ (.A(_3162_),
    .B(_3164_),
    .X(_3165_));
 sky130_fd_sc_hd__nand2_1 _7989_ (.A(_3162_),
    .B(_3164_),
    .Y(_3166_));
 sky130_fd_sc_hd__xor2_1 _7990_ (.A(_3149_),
    .B(_3151_),
    .X(_3167_));
 sky130_fd_sc_hd__xnor2_1 _7991_ (.A(_3153_),
    .B(_3167_),
    .Y(_3169_));
 sky130_fd_sc_hd__a21o_1 _7992_ (.A1(net13),
    .A2(_1760_),
    .B1(_3169_),
    .X(_3170_));
 sky130_fd_sc_hd__or3b_1 _7993_ (.A(_0000_),
    .B(_1771_),
    .C_N(_3169_),
    .X(_3171_));
 sky130_fd_sc_hd__and2b_1 _7994_ (.A_N(_3005_),
    .B(_3006_),
    .X(_3172_));
 sky130_fd_sc_hd__xor2_1 _7995_ (.A(_3148_),
    .B(_3172_),
    .X(_3173_));
 sky130_fd_sc_hd__xor2_1 _7996_ (.A(_3141_),
    .B(_3143_),
    .X(_3174_));
 sky130_fd_sc_hd__xnor2_1 _7997_ (.A(_3145_),
    .B(_3174_),
    .Y(_3175_));
 sky130_fd_sc_hd__a21o_1 _7998_ (.A1(net10),
    .A2(_1760_),
    .B1(_3175_),
    .X(_3176_));
 sky130_fd_sc_hd__nand3_1 _7999_ (.A(net10),
    .B(_1760_),
    .C(_3175_),
    .Y(_3177_));
 sky130_fd_sc_hd__nor2_1 _8000_ (.A(_3011_),
    .B(_3013_),
    .Y(_3178_));
 sky130_fd_sc_hd__xnor2_1 _8001_ (.A(_3140_),
    .B(_3178_),
    .Y(_3180_));
 sky130_fd_sc_hd__nand2_1 _8002_ (.A(net8),
    .B(_1760_),
    .Y(_3181_));
 sky130_fd_sc_hd__xor2_1 _8003_ (.A(_3133_),
    .B(_3136_),
    .X(_3182_));
 sky130_fd_sc_hd__xnor2_1 _8004_ (.A(_3138_),
    .B(_3182_),
    .Y(_3183_));
 sky130_fd_sc_hd__nand2_1 _8005_ (.A(_3181_),
    .B(_3183_),
    .Y(_3184_));
 sky130_fd_sc_hd__or2_1 _8006_ (.A(_3181_),
    .B(_3183_),
    .X(_3185_));
 sky130_fd_sc_hd__nor2_1 _8007_ (.A(_3019_),
    .B(_3021_),
    .Y(_3186_));
 sky130_fd_sc_hd__xnor2_1 _8008_ (.A(_3131_),
    .B(_3186_),
    .Y(_3187_));
 sky130_fd_sc_hd__xor2_1 _8009_ (.A(_3125_),
    .B(_3127_),
    .X(_3188_));
 sky130_fd_sc_hd__xnor2_1 _8010_ (.A(_3129_),
    .B(_3188_),
    .Y(_3189_));
 sky130_fd_sc_hd__nor2_1 _8011_ (.A(_3026_),
    .B(_3028_),
    .Y(_3191_));
 sky130_fd_sc_hd__xnor2_1 _8012_ (.A(_3123_),
    .B(_3191_),
    .Y(_3192_));
 sky130_fd_sc_hd__xnor2_1 _8013_ (.A(_3117_),
    .B(_3119_),
    .Y(_3193_));
 sky130_fd_sc_hd__xnor2_1 _8014_ (.A(_3121_),
    .B(_3193_),
    .Y(_3194_));
 sky130_fd_sc_hd__xor2_1 _8015_ (.A(_3029_),
    .B(_3032_),
    .X(_3195_));
 sky130_fd_sc_hd__xnor2_1 _8016_ (.A(_3115_),
    .B(_3195_),
    .Y(_3196_));
 sky130_fd_sc_hd__xor2_1 _8017_ (.A(_3108_),
    .B(_3110_),
    .X(_3197_));
 sky130_fd_sc_hd__xnor2_1 _8018_ (.A(_3112_),
    .B(_3197_),
    .Y(_3198_));
 sky130_fd_sc_hd__nand2b_1 _8019_ (.A_N(_3040_),
    .B(_3041_),
    .Y(_3199_));
 sky130_fd_sc_hd__xnor2_1 _8020_ (.A(_3107_),
    .B(_3199_),
    .Y(_3200_));
 sky130_fd_sc_hd__xor2_1 _8021_ (.A(_3100_),
    .B(_3103_),
    .X(_3202_));
 sky130_fd_sc_hd__xnor2_1 _8022_ (.A(_3105_),
    .B(_3202_),
    .Y(_3203_));
 sky130_fd_sc_hd__nand2b_1 _8023_ (.A_N(_3045_),
    .B(_3046_),
    .Y(_3204_));
 sky130_fd_sc_hd__xor2_1 _8024_ (.A(_3099_),
    .B(_3204_),
    .X(_3205_));
 sky130_fd_sc_hd__xor2_1 _8025_ (.A(_3093_),
    .B(_3095_),
    .X(_3206_));
 sky130_fd_sc_hd__xor2_1 _8026_ (.A(_3097_),
    .B(_3206_),
    .X(_3207_));
 sky130_fd_sc_hd__xnor2_1 _8027_ (.A(_3048_),
    .B(_3051_),
    .Y(_3208_));
 sky130_fd_sc_hd__xor2_1 _8028_ (.A(_3092_),
    .B(_3208_),
    .X(_3209_));
 sky130_fd_sc_hd__xor2_1 _8029_ (.A(_3085_),
    .B(_3087_),
    .X(_3210_));
 sky130_fd_sc_hd__xor2_2 _8030_ (.A(_3089_),
    .B(_3210_),
    .X(_3211_));
 sky130_fd_sc_hd__nor2_1 _8031_ (.A(_3057_),
    .B(_3060_),
    .Y(_3213_));
 sky130_fd_sc_hd__xnor2_2 _8032_ (.A(_3084_),
    .B(_3213_),
    .Y(_3214_));
 sky130_fd_sc_hd__xor2_1 _8033_ (.A(_3061_),
    .B(_3063_),
    .X(_3215_));
 sky130_fd_sc_hd__xnor2_1 _8034_ (.A(_3076_),
    .B(_3215_),
    .Y(_3216_));
 sky130_fd_sc_hd__a21bo_1 _8035_ (.A1(net12),
    .A2(_1760_),
    .B1_N(_3216_),
    .X(_3217_));
 sky130_fd_sc_hd__inv_2 _8036_ (.A(_3217_),
    .Y(_3218_));
 sky130_fd_sc_hd__nor3b_1 _8037_ (.A(_1771_),
    .B(_3216_),
    .C_N(net12),
    .Y(_3219_));
 sky130_fd_sc_hd__nor2_1 _8038_ (.A(_3070_),
    .B(_3072_),
    .Y(_3220_));
 sky130_fd_sc_hd__xnor2_1 _8039_ (.A(_3075_),
    .B(_3220_),
    .Y(_3221_));
 sky130_fd_sc_hd__and3b_1 _8040_ (.A_N(_3221_),
    .B(net1),
    .C(_1760_),
    .X(_3222_));
 sky130_fd_sc_hd__a21o_1 _8041_ (.A1(_3217_),
    .A2(_3222_),
    .B1(_3219_),
    .X(_3224_));
 sky130_fd_sc_hd__xor2_1 _8042_ (.A(_3077_),
    .B(_3079_),
    .X(_3225_));
 sky130_fd_sc_hd__xnor2_1 _8043_ (.A(_3082_),
    .B(_3225_),
    .Y(_3226_));
 sky130_fd_sc_hd__or2_2 _8044_ (.A(_3224_),
    .B(_3226_),
    .X(_3227_));
 sky130_fd_sc_hd__inv_2 _8045_ (.A(_3227_),
    .Y(_3228_));
 sky130_fd_sc_hd__and2_1 _8046_ (.A(_3224_),
    .B(_3226_),
    .X(_3229_));
 sky130_fd_sc_hd__and2_1 _8047_ (.A(net23),
    .B(_1760_),
    .X(_3230_));
 sky130_fd_sc_hd__a21o_1 _8048_ (.A1(_3224_),
    .A2(_3226_),
    .B1(_3230_),
    .X(_3231_));
 sky130_fd_sc_hd__a21oi_2 _8049_ (.A1(_3227_),
    .A2(_3231_),
    .B1(_3214_),
    .Y(_3232_));
 sky130_fd_sc_hd__and3_1 _8050_ (.A(_3214_),
    .B(_3227_),
    .C(_3231_),
    .X(_3233_));
 sky130_fd_sc_hd__nand2_1 _8051_ (.A(net26),
    .B(_1760_),
    .Y(_3235_));
 sky130_fd_sc_hd__inv_2 _8052_ (.A(_3235_),
    .Y(_3236_));
 sky130_fd_sc_hd__a31oi_2 _8053_ (.A1(_3214_),
    .A2(_3227_),
    .A3(_3231_),
    .B1(_3236_),
    .Y(_3237_));
 sky130_fd_sc_hd__o21ai_2 _8054_ (.A1(_3232_),
    .A2(_3237_),
    .B1(_3211_),
    .Y(_3238_));
 sky130_fd_sc_hd__or3_1 _8055_ (.A(_3211_),
    .B(_3232_),
    .C(_3237_),
    .X(_3239_));
 sky130_fd_sc_hd__nor2_1 _8056_ (.A(_4187_),
    .B(_1771_),
    .Y(_3240_));
 sky130_fd_sc_hd__o32ai_2 _8057_ (.A1(_3211_),
    .A2(_3232_),
    .A3(_3237_),
    .B1(_1771_),
    .B2(_4187_),
    .Y(_3241_));
 sky130_fd_sc_hd__a21o_1 _8058_ (.A1(_3238_),
    .A2(_3241_),
    .B1(_3209_),
    .X(_3242_));
 sky130_fd_sc_hd__nand3_1 _8059_ (.A(_3209_),
    .B(_3238_),
    .C(_3241_),
    .Y(_3243_));
 sky130_fd_sc_hd__nand2_1 _8060_ (.A(net28),
    .B(_1760_),
    .Y(_3244_));
 sky130_fd_sc_hd__a32o_1 _8061_ (.A1(_3209_),
    .A2(_3238_),
    .A3(_3241_),
    .B1(_1760_),
    .B2(net28),
    .X(_3246_));
 sky130_fd_sc_hd__a21o_1 _8062_ (.A1(_3242_),
    .A2(_3246_),
    .B1(_3207_),
    .X(_3247_));
 sky130_fd_sc_hd__nand3_1 _8063_ (.A(_3207_),
    .B(_3242_),
    .C(_3246_),
    .Y(_3248_));
 sky130_fd_sc_hd__and2_1 _8064_ (.A(net29),
    .B(_1760_),
    .X(_3249_));
 sky130_fd_sc_hd__a31o_1 _8065_ (.A1(_3207_),
    .A2(_3242_),
    .A3(_3246_),
    .B1(_3249_),
    .X(_3250_));
 sky130_fd_sc_hd__a21o_1 _8066_ (.A1(_3247_),
    .A2(_3250_),
    .B1(_3205_),
    .X(_3251_));
 sky130_fd_sc_hd__nand3_1 _8067_ (.A(_3205_),
    .B(_3247_),
    .C(_3250_),
    .Y(_3252_));
 sky130_fd_sc_hd__nand2_1 _8068_ (.A(net30),
    .B(_1760_),
    .Y(_3253_));
 sky130_fd_sc_hd__inv_2 _8069_ (.A(_3253_),
    .Y(_3254_));
 sky130_fd_sc_hd__a31o_1 _8070_ (.A1(_3205_),
    .A2(_3247_),
    .A3(_3250_),
    .B1(_3254_),
    .X(_3255_));
 sky130_fd_sc_hd__a21oi_1 _8071_ (.A1(_3251_),
    .A2(_3255_),
    .B1(_3203_),
    .Y(_3257_));
 sky130_fd_sc_hd__a21o_1 _8072_ (.A1(_3251_),
    .A2(_3255_),
    .B1(_3203_),
    .X(_3258_));
 sky130_fd_sc_hd__and3_1 _8073_ (.A(_3203_),
    .B(_3251_),
    .C(_3255_),
    .X(_3259_));
 sky130_fd_sc_hd__nand2_1 _8074_ (.A(net31),
    .B(_1760_),
    .Y(_3260_));
 sky130_fd_sc_hd__a32o_1 _8075_ (.A1(_3203_),
    .A2(_3251_),
    .A3(_3255_),
    .B1(_1760_),
    .B2(net31),
    .X(_3261_));
 sky130_fd_sc_hd__a21o_1 _8076_ (.A1(_3258_),
    .A2(_3261_),
    .B1(_3200_),
    .X(_3262_));
 sky130_fd_sc_hd__nand3_1 _8077_ (.A(_3200_),
    .B(_3258_),
    .C(_3261_),
    .Y(_3263_));
 sky130_fd_sc_hd__nand2_1 _8078_ (.A(net32),
    .B(_1760_),
    .Y(_3264_));
 sky130_fd_sc_hd__a32o_1 _8079_ (.A1(_3200_),
    .A2(_3258_),
    .A3(_3261_),
    .B1(_1760_),
    .B2(net32),
    .X(_3265_));
 sky130_fd_sc_hd__a21o_1 _8080_ (.A1(_3262_),
    .A2(_3265_),
    .B1(_3198_),
    .X(_3266_));
 sky130_fd_sc_hd__nand3_1 _8081_ (.A(_3198_),
    .B(_3262_),
    .C(_3265_),
    .Y(_3268_));
 sky130_fd_sc_hd__and2_1 _8082_ (.A(net2),
    .B(_1760_),
    .X(_3269_));
 sky130_fd_sc_hd__a31o_1 _8083_ (.A1(_3198_),
    .A2(_3262_),
    .A3(_3265_),
    .B1(_3269_),
    .X(_3270_));
 sky130_fd_sc_hd__a21o_1 _8084_ (.A1(_3266_),
    .A2(_3270_),
    .B1(_3196_),
    .X(_3271_));
 sky130_fd_sc_hd__nand3_1 _8085_ (.A(_3196_),
    .B(_3266_),
    .C(_3270_),
    .Y(_3272_));
 sky130_fd_sc_hd__nand2_1 _8086_ (.A(net3),
    .B(_1760_),
    .Y(_3273_));
 sky130_fd_sc_hd__a32o_1 _8087_ (.A1(_3196_),
    .A2(_3266_),
    .A3(_3270_),
    .B1(_1760_),
    .B2(net3),
    .X(_3274_));
 sky130_fd_sc_hd__a21o_1 _8088_ (.A1(_3271_),
    .A2(_3274_),
    .B1(_3194_),
    .X(_3275_));
 sky130_fd_sc_hd__nand3_1 _8089_ (.A(_3194_),
    .B(_3271_),
    .C(_3274_),
    .Y(_3276_));
 sky130_fd_sc_hd__and2_1 _8090_ (.A(net4),
    .B(_1760_),
    .X(_3277_));
 sky130_fd_sc_hd__a31o_1 _8091_ (.A1(_3194_),
    .A2(_3271_),
    .A3(_3274_),
    .B1(_3277_),
    .X(_3279_));
 sky130_fd_sc_hd__a21o_1 _8092_ (.A1(_3275_),
    .A2(_3279_),
    .B1(_3192_),
    .X(_3280_));
 sky130_fd_sc_hd__nand3_1 _8093_ (.A(_3192_),
    .B(_3275_),
    .C(_3279_),
    .Y(_3281_));
 sky130_fd_sc_hd__nand2_1 _8094_ (.A(net5),
    .B(_1760_),
    .Y(_3282_));
 sky130_fd_sc_hd__a32o_1 _8095_ (.A1(_3192_),
    .A2(_3275_),
    .A3(_3279_),
    .B1(_1760_),
    .B2(net5),
    .X(_3283_));
 sky130_fd_sc_hd__a21o_1 _8096_ (.A1(_3280_),
    .A2(_3283_),
    .B1(_3189_),
    .X(_3284_));
 sky130_fd_sc_hd__nand3_1 _8097_ (.A(_3189_),
    .B(_3280_),
    .C(_3283_),
    .Y(_3285_));
 sky130_fd_sc_hd__nand2_1 _8098_ (.A(net6),
    .B(_1760_),
    .Y(_3286_));
 sky130_fd_sc_hd__a32o_1 _8099_ (.A1(_3189_),
    .A2(_3280_),
    .A3(_3283_),
    .B1(_1760_),
    .B2(net6),
    .X(_3287_));
 sky130_fd_sc_hd__a21o_1 _8100_ (.A1(_3284_),
    .A2(_3287_),
    .B1(_3187_),
    .X(_3288_));
 sky130_fd_sc_hd__nand3_1 _8101_ (.A(_3187_),
    .B(_3284_),
    .C(_3287_),
    .Y(_3290_));
 sky130_fd_sc_hd__nand2_1 _8102_ (.A(net7),
    .B(_1760_),
    .Y(_3291_));
 sky130_fd_sc_hd__a32o_1 _8103_ (.A1(_3187_),
    .A2(_3284_),
    .A3(_3287_),
    .B1(_1760_),
    .B2(net7),
    .X(_3292_));
 sky130_fd_sc_hd__and2_1 _8104_ (.A(_3288_),
    .B(_3292_),
    .X(_3293_));
 sky130_fd_sc_hd__a2bb2o_1 _8105_ (.A1_N(_3181_),
    .A2_N(_3183_),
    .B1(_3288_),
    .B2(_3292_),
    .X(_3294_));
 sky130_fd_sc_hd__a21o_1 _8106_ (.A1(_3184_),
    .A2(_3294_),
    .B1(_3180_),
    .X(_3295_));
 sky130_fd_sc_hd__nand3_1 _8107_ (.A(_3180_),
    .B(_3184_),
    .C(_3294_),
    .Y(_3296_));
 sky130_fd_sc_hd__nand2_1 _8108_ (.A(net9),
    .B(_1760_),
    .Y(_3297_));
 sky130_fd_sc_hd__inv_2 _8109_ (.A(_3297_),
    .Y(_3298_));
 sky130_fd_sc_hd__a31o_1 _8110_ (.A1(_3180_),
    .A2(_3184_),
    .A3(_3294_),
    .B1(_3298_),
    .X(_3299_));
 sky130_fd_sc_hd__nand2_1 _8111_ (.A(_3295_),
    .B(_3299_),
    .Y(_3301_));
 sky130_fd_sc_hd__a32o_1 _8112_ (.A1(net10),
    .A2(_1760_),
    .A3(_3175_),
    .B1(_3295_),
    .B2(_3299_),
    .X(_3302_));
 sky130_fd_sc_hd__a21o_1 _8113_ (.A1(_3176_),
    .A2(_3302_),
    .B1(_3173_),
    .X(_3303_));
 sky130_fd_sc_hd__nand3_1 _8114_ (.A(_3173_),
    .B(_3176_),
    .C(_3302_),
    .Y(_3304_));
 sky130_fd_sc_hd__nand2_1 _8115_ (.A(net11),
    .B(_1760_),
    .Y(_3305_));
 sky130_fd_sc_hd__a32o_1 _8116_ (.A1(_3173_),
    .A2(_3176_),
    .A3(_3302_),
    .B1(_1760_),
    .B2(net11),
    .X(_3306_));
 sky130_fd_sc_hd__nand2_1 _8117_ (.A(_3303_),
    .B(_3306_),
    .Y(_3307_));
 sky130_fd_sc_hd__a32o_1 _8118_ (.A1(net13),
    .A2(_1760_),
    .A3(_3169_),
    .B1(_3303_),
    .B2(_3306_),
    .X(_3308_));
 sky130_fd_sc_hd__and2b_1 _8119_ (.A_N(_3000_),
    .B(_3001_),
    .X(_3309_));
 sky130_fd_sc_hd__xor2_1 _8120_ (.A(_3155_),
    .B(_3309_),
    .X(_3310_));
 sky130_fd_sc_hd__a21o_1 _8121_ (.A1(_3170_),
    .A2(_3308_),
    .B1(_3310_),
    .X(_3312_));
 sky130_fd_sc_hd__nand3_1 _8122_ (.A(_3170_),
    .B(_3308_),
    .C(_3310_),
    .Y(_3313_));
 sky130_fd_sc_hd__nand2_1 _8123_ (.A(net14),
    .B(_1760_),
    .Y(_3314_));
 sky130_fd_sc_hd__inv_2 _8124_ (.A(_3314_),
    .Y(_3315_));
 sky130_fd_sc_hd__a31o_1 _8125_ (.A1(_3170_),
    .A2(_3308_),
    .A3(_3310_),
    .B1(_3315_),
    .X(_3316_));
 sky130_fd_sc_hd__and2_1 _8126_ (.A(_3312_),
    .B(_3316_),
    .X(_3317_));
 sky130_fd_sc_hd__a22o_1 _8127_ (.A1(_3162_),
    .A2(_3164_),
    .B1(_3312_),
    .B2(_3316_),
    .X(_3318_));
 sky130_fd_sc_hd__nand2_1 _8128_ (.A(_3165_),
    .B(_3318_),
    .Y(_3319_));
 sky130_fd_sc_hd__a32o_4 _8129_ (.A1(_3160_),
    .A2(_3165_),
    .A3(_3318_),
    .B1(_3159_),
    .B2(_1760_),
    .X(_3320_));
 sky130_fd_sc_hd__and2_1 _8130_ (.A(_0638_),
    .B(_3972_),
    .X(_3321_));
 sky130_fd_sc_hd__xor2_2 _8131_ (.A(_3960_),
    .B(_3961_),
    .X(_3323_));
 sky130_fd_sc_hd__xnor2_1 _8132_ (.A(_3957_),
    .B(_3962_),
    .Y(_3324_));
 sky130_fd_sc_hd__and4_2 _8133_ (.A(_3320_),
    .B(_3321_),
    .C(_3323_),
    .D(_3324_),
    .X(_3325_));
 sky130_fd_sc_hd__nor2_1 _8134_ (.A(_3954_),
    .B(_3966_),
    .Y(_3326_));
 sky130_fd_sc_hd__and3_1 _8135_ (.A(_3970_),
    .B(_3325_),
    .C(_3326_),
    .X(_3327_));
 sky130_fd_sc_hd__a21oi_1 _8136_ (.A1(_3325_),
    .A2(_3326_),
    .B1(_3970_),
    .Y(_3328_));
 sky130_fd_sc_hd__and2_1 _8137_ (.A(_3963_),
    .B(_3966_),
    .X(_3329_));
 sky130_fd_sc_hd__nor2_1 _8138_ (.A(_3967_),
    .B(_3329_),
    .Y(_3330_));
 sky130_fd_sc_hd__nor2_1 _8139_ (.A(_3964_),
    .B(_3967_),
    .Y(_3331_));
 sky130_fd_sc_hd__xnor2_1 _8140_ (.A(_3954_),
    .B(_3331_),
    .Y(_3332_));
 sky130_fd_sc_hd__a21oi_1 _8141_ (.A1(_3325_),
    .A2(_3330_),
    .B1(_3332_),
    .Y(_3334_));
 sky130_fd_sc_hd__xnor2_1 _8142_ (.A(_0649_),
    .B(_3320_),
    .Y(_3335_));
 sky130_fd_sc_hd__a221o_1 _8143_ (.A1(net22),
    .A2(net54),
    .B1(_3950_),
    .B2(_3969_),
    .C1(_3948_),
    .X(_3336_));
 sky130_fd_sc_hd__xor2_1 _8144_ (.A(_0836_),
    .B(_3336_),
    .X(_3337_));
 sky130_fd_sc_hd__and4_1 _8145_ (.A(_3960_),
    .B(_3972_),
    .C(_3330_),
    .D(_3337_),
    .X(_3338_));
 sky130_fd_sc_hd__nand2_1 _8146_ (.A(_3335_),
    .B(_3338_),
    .Y(_3339_));
 sky130_fd_sc_hd__a31o_1 _8147_ (.A1(_3320_),
    .A2(_3321_),
    .A3(_3323_),
    .B1(_3324_),
    .X(_3340_));
 sky130_fd_sc_hd__or3b_1 _8148_ (.A(_3325_),
    .B(_3332_),
    .C_N(_3340_),
    .X(_3341_));
 sky130_fd_sc_hd__or4_4 _8149_ (.A(_3327_),
    .B(_3328_),
    .C(_3339_),
    .D(_3341_),
    .X(_3342_));
 sky130_fd_sc_hd__nand2_4 _8150_ (.A(_3944_),
    .B(_3945_),
    .Y(_3343_));
 sky130_fd_sc_hd__nor2_1 _8151_ (.A(_0462_),
    .B(_3343_),
    .Y(_3345_));
 sky130_fd_sc_hd__and3_4 _8152_ (.A(_3947_),
    .B(_3342_),
    .C(_3345_),
    .X(_3346_));
 sky130_fd_sc_hd__nor2_1 _8153_ (.A(_3218_),
    .B(_3219_),
    .Y(_3347_));
 sky130_fd_sc_hd__xor2_1 _8154_ (.A(_3222_),
    .B(_3347_),
    .X(_3348_));
 sky130_fd_sc_hd__or2_1 _8155_ (.A(net24),
    .B(net56),
    .X(_3349_));
 sky130_fd_sc_hd__nor2_2 _8156_ (.A(_3336_),
    .B(_3349_),
    .Y(_3350_));
 sky130_fd_sc_hd__or2_4 _8157_ (.A(_3336_),
    .B(_3349_),
    .X(_3351_));
 sky130_fd_sc_hd__o21a_1 _8158_ (.A1(_4198_),
    .A2(_1771_),
    .B1(_3221_),
    .X(_3352_));
 sky130_fd_sc_hd__nand2_1 _8159_ (.A(_3320_),
    .B(_3348_),
    .Y(_3353_));
 sky130_fd_sc_hd__o31ai_2 _8160_ (.A1(_3222_),
    .A2(_3320_),
    .A3(_3352_),
    .B1(_3353_),
    .Y(_3354_));
 sky130_fd_sc_hd__a31o_1 _8161_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3354_),
    .B1(_3943_),
    .X(net66));
 sky130_fd_sc_hd__nand2b_1 _8162_ (.A_N(_3900_),
    .B(_3902_),
    .Y(_3356_));
 sky130_fd_sc_hd__nand2_1 _8163_ (.A(_3903_),
    .B(_3356_),
    .Y(_3357_));
 sky130_fd_sc_hd__nor3_1 _8164_ (.A(_3932_),
    .B(_3934_),
    .C(_3936_),
    .Y(_3358_));
 sky130_fd_sc_hd__a21bo_1 _8165_ (.A1(_3753_),
    .A2(_3938_),
    .B1_N(_1122_),
    .X(_3359_));
 sky130_fd_sc_hd__a211oi_1 _8166_ (.A1(_3932_),
    .A2(_3357_),
    .B1(_3358_),
    .C1(_3359_),
    .Y(_3360_));
 sky130_fd_sc_hd__nor2_1 _8167_ (.A(_3228_),
    .B(_3229_),
    .Y(_3361_));
 sky130_fd_sc_hd__xnor2_1 _8168_ (.A(_3230_),
    .B(_3361_),
    .Y(_3362_));
 sky130_fd_sc_hd__inv_2 _8169_ (.A(_3362_),
    .Y(_3363_));
 sky130_fd_sc_hd__mux2_1 _8170_ (.A0(_3348_),
    .A1(_3363_),
    .S(_3320_),
    .X(_3364_));
 sky130_fd_sc_hd__a31o_1 _8171_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3364_),
    .B1(_3360_),
    .X(net77));
 sky130_fd_sc_hd__nor2_1 _8172_ (.A(_3232_),
    .B(_3233_),
    .Y(_3366_));
 sky130_fd_sc_hd__xnor2_1 _8173_ (.A(_3236_),
    .B(_3366_),
    .Y(_3367_));
 sky130_fd_sc_hd__nand2_1 _8174_ (.A(_3320_),
    .B(_3367_),
    .Y(_3368_));
 sky130_fd_sc_hd__o211a_1 _8175_ (.A1(_3320_),
    .A2(_3363_),
    .B1(_3368_),
    .C1(_3351_),
    .X(_3369_));
 sky130_fd_sc_hd__and3_1 _8176_ (.A(_3820_),
    .B(_3823_),
    .C(_3926_),
    .X(_3370_));
 sky130_fd_sc_hd__or2_1 _8177_ (.A(_3927_),
    .B(_3370_),
    .X(_3371_));
 sky130_fd_sc_hd__or3_1 _8178_ (.A(_3825_),
    .B(_3828_),
    .C(_3925_),
    .X(_3372_));
 sky130_fd_sc_hd__nand2_1 _8179_ (.A(_3926_),
    .B(_3372_),
    .Y(_3373_));
 sky130_fd_sc_hd__xnor2_1 _8180_ (.A(_3830_),
    .B(_3924_),
    .Y(_3374_));
 sky130_fd_sc_hd__and3_1 _8181_ (.A(_3833_),
    .B(_3836_),
    .C(_3922_),
    .X(_3376_));
 sky130_fd_sc_hd__or2_1 _8182_ (.A(_3923_),
    .B(_3376_),
    .X(_3377_));
 sky130_fd_sc_hd__or3_1 _8183_ (.A(_3838_),
    .B(_3841_),
    .C(_3921_),
    .X(_3378_));
 sky130_fd_sc_hd__nand2_1 _8184_ (.A(_3922_),
    .B(_3378_),
    .Y(_3379_));
 sky130_fd_sc_hd__nor3_1 _8185_ (.A(_3842_),
    .B(_3845_),
    .C(_3920_),
    .Y(_3380_));
 sky130_fd_sc_hd__or2_1 _8186_ (.A(_3921_),
    .B(_3380_),
    .X(_3381_));
 sky130_fd_sc_hd__and3_1 _8187_ (.A(_3846_),
    .B(_3849_),
    .C(_3919_),
    .X(_3382_));
 sky130_fd_sc_hd__or2_1 _8188_ (.A(_3920_),
    .B(_3382_),
    .X(_3383_));
 sky130_fd_sc_hd__nand3_1 _8189_ (.A(_3850_),
    .B(_3853_),
    .C(_3918_),
    .Y(_3384_));
 sky130_fd_sc_hd__nand2_1 _8190_ (.A(_3919_),
    .B(_3384_),
    .Y(_3385_));
 sky130_fd_sc_hd__or3_1 _8191_ (.A(_3855_),
    .B(_3858_),
    .C(_3917_),
    .X(_3387_));
 sky130_fd_sc_hd__nand2_1 _8192_ (.A(_3918_),
    .B(_3387_),
    .Y(_3388_));
 sky130_fd_sc_hd__xnor2_2 _8193_ (.A(_3860_),
    .B(_3916_),
    .Y(_3389_));
 sky130_fd_sc_hd__or3_1 _8194_ (.A(_3864_),
    .B(_3867_),
    .C(_3914_),
    .X(_3390_));
 sky130_fd_sc_hd__nand2_1 _8195_ (.A(_3915_),
    .B(_3390_),
    .Y(_3391_));
 sky130_fd_sc_hd__xnor2_1 _8196_ (.A(_3869_),
    .B(_3913_),
    .Y(_3392_));
 sky130_fd_sc_hd__and3_1 _8197_ (.A(_3872_),
    .B(_3875_),
    .C(_3911_),
    .X(_3393_));
 sky130_fd_sc_hd__nor2_1 _8198_ (.A(_3912_),
    .B(_3393_),
    .Y(_3394_));
 sky130_fd_sc_hd__xnor2_2 _8199_ (.A(_3876_),
    .B(_3910_),
    .Y(_3395_));
 sky130_fd_sc_hd__or3_1 _8200_ (.A(_3880_),
    .B(_3883_),
    .C(_3908_),
    .X(_3396_));
 sky130_fd_sc_hd__and2_1 _8201_ (.A(_3909_),
    .B(_3396_),
    .X(_3398_));
 sky130_fd_sc_hd__xnor2_1 _8202_ (.A(_3884_),
    .B(_3907_),
    .Y(_3399_));
 sky130_fd_sc_hd__and3_1 _8203_ (.A(_3887_),
    .B(_3890_),
    .C(_3905_),
    .X(_3400_));
 sky130_fd_sc_hd__nor2_1 _8204_ (.A(_3906_),
    .B(_3400_),
    .Y(_3401_));
 sky130_fd_sc_hd__nand3_1 _8205_ (.A(_3891_),
    .B(_3894_),
    .C(_3904_),
    .Y(_3402_));
 sky130_fd_sc_hd__nand2_1 _8206_ (.A(_3905_),
    .B(_3402_),
    .Y(_3403_));
 sky130_fd_sc_hd__inv_2 _8207_ (.A(_3403_),
    .Y(_3404_));
 sky130_fd_sc_hd__nand3_1 _8208_ (.A(_3896_),
    .B(_3899_),
    .C(_3903_),
    .Y(_3405_));
 sky130_fd_sc_hd__and2_1 _8209_ (.A(_3904_),
    .B(_3405_),
    .X(_3406_));
 sky130_fd_sc_hd__nand2_1 _8210_ (.A(_3753_),
    .B(_3357_),
    .Y(_3407_));
 sky130_fd_sc_hd__or4_1 _8211_ (.A(_3401_),
    .B(_3404_),
    .C(_3406_),
    .D(_3407_),
    .X(_3409_));
 sky130_fd_sc_hd__or4_1 _8212_ (.A(_3395_),
    .B(_3398_),
    .C(_3399_),
    .D(_3409_),
    .X(_3410_));
 sky130_fd_sc_hd__or4b_1 _8213_ (.A(_3392_),
    .B(_3410_),
    .C(_3394_),
    .D_N(_3391_),
    .X(_3411_));
 sky130_fd_sc_hd__and4b_1 _8214_ (.A_N(_3411_),
    .B(_3389_),
    .C(_3388_),
    .D(_3385_),
    .X(_3412_));
 sky130_fd_sc_hd__and4_1 _8215_ (.A(_3379_),
    .B(_3381_),
    .C(_3383_),
    .D(_3412_),
    .X(_3413_));
 sky130_fd_sc_hd__and4_1 _8216_ (.A(_3373_),
    .B(_3374_),
    .C(_3377_),
    .D(_3413_),
    .X(_3414_));
 sky130_fd_sc_hd__xnor2_2 _8217_ (.A(_3817_),
    .B(_3928_),
    .Y(_3415_));
 sky130_fd_sc_hd__and4_2 _8218_ (.A(_3358_),
    .B(_3371_),
    .C(_3414_),
    .D(_3415_),
    .X(_3416_));
 sky130_fd_sc_hd__and2b_4 _8219_ (.A_N(_3416_),
    .B(_1122_),
    .X(_3417_));
 sky130_fd_sc_hd__nand2_1 _8220_ (.A(_3938_),
    .B(_3357_),
    .Y(_3418_));
 sky130_fd_sc_hd__nand2_1 _8221_ (.A(_3753_),
    .B(_3937_),
    .Y(_3420_));
 sky130_fd_sc_hd__mux2_1 _8222_ (.A0(_3420_),
    .A1(_3406_),
    .S(_3932_),
    .X(_3421_));
 sky130_fd_sc_hd__a32o_1 _8223_ (.A1(_3417_),
    .A2(_3418_),
    .A3(_3421_),
    .B1(_3369_),
    .B2(_3346_),
    .X(net88));
 sky130_fd_sc_hd__nor2_1 _8224_ (.A(_3320_),
    .B(_3367_),
    .Y(_3422_));
 sky130_fd_sc_hd__nand2_1 _8225_ (.A(_3238_),
    .B(_3239_),
    .Y(_3423_));
 sky130_fd_sc_hd__xnor2_1 _8226_ (.A(_3240_),
    .B(_3423_),
    .Y(_3424_));
 sky130_fd_sc_hd__a21o_1 _8227_ (.A1(_3320_),
    .A2(_3424_),
    .B1(_3422_),
    .X(_3425_));
 sky130_fd_sc_hd__nand2_1 _8228_ (.A(_3937_),
    .B(_3357_),
    .Y(_3426_));
 sky130_fd_sc_hd__mux2_1 _8229_ (.A0(_3426_),
    .A1(_3404_),
    .S(_3932_),
    .X(_3427_));
 sky130_fd_sc_hd__o211a_1 _8230_ (.A1(_3939_),
    .A2(_3406_),
    .B1(_3417_),
    .C1(_3427_),
    .X(_3428_));
 sky130_fd_sc_hd__a31o_1 _8231_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3425_),
    .B1(_3428_),
    .X(net91));
 sky130_fd_sc_hd__nand2_1 _8232_ (.A(_3242_),
    .B(_3243_),
    .Y(_3430_));
 sky130_fd_sc_hd__xor2_1 _8233_ (.A(_3244_),
    .B(_3430_),
    .X(_3431_));
 sky130_fd_sc_hd__mux2_1 _8234_ (.A0(_3424_),
    .A1(_3431_),
    .S(_3320_),
    .X(_3432_));
 sky130_fd_sc_hd__nand2_1 _8235_ (.A(_3938_),
    .B(_3403_),
    .Y(_3433_));
 sky130_fd_sc_hd__or3_1 _8236_ (.A(_3932_),
    .B(_3936_),
    .C(_3406_),
    .X(_3434_));
 sky130_fd_sc_hd__o2111a_1 _8237_ (.A1(_3933_),
    .A2(_3401_),
    .B1(_3417_),
    .C1(_3433_),
    .D1(_3434_),
    .X(_3435_));
 sky130_fd_sc_hd__a31o_1 _8238_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3432_),
    .B1(_3435_),
    .X(net92));
 sky130_fd_sc_hd__nand2_1 _8239_ (.A(_3247_),
    .B(_3248_),
    .Y(_3436_));
 sky130_fd_sc_hd__xor2_1 _8240_ (.A(_3249_),
    .B(_3436_),
    .X(_3437_));
 sky130_fd_sc_hd__inv_2 _8241_ (.A(_3437_),
    .Y(_3439_));
 sky130_fd_sc_hd__mux2_1 _8242_ (.A0(_3431_),
    .A1(_3439_),
    .S(_3320_),
    .X(_3440_));
 sky130_fd_sc_hd__nand2_1 _8243_ (.A(_3937_),
    .B(_3403_),
    .Y(_3441_));
 sky130_fd_sc_hd__mux2_1 _8244_ (.A0(_3441_),
    .A1(_3399_),
    .S(_3932_),
    .X(_3442_));
 sky130_fd_sc_hd__o211a_1 _8245_ (.A1(_3939_),
    .A2(_3401_),
    .B1(_3417_),
    .C1(_3442_),
    .X(_3443_));
 sky130_fd_sc_hd__a31o_1 _8246_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3440_),
    .B1(_3443_),
    .X(net93));
 sky130_fd_sc_hd__nand2_1 _8247_ (.A(_3251_),
    .B(_3252_),
    .Y(_3444_));
 sky130_fd_sc_hd__xnor2_1 _8248_ (.A(_3254_),
    .B(_3444_),
    .Y(_3445_));
 sky130_fd_sc_hd__mux2_1 _8249_ (.A0(_3439_),
    .A1(_3445_),
    .S(_3320_),
    .X(_3446_));
 sky130_fd_sc_hd__or2_1 _8250_ (.A(_3939_),
    .B(_3399_),
    .X(_3447_));
 sky130_fd_sc_hd__or3_1 _8251_ (.A(_3932_),
    .B(_3936_),
    .C(_3401_),
    .X(_3449_));
 sky130_fd_sc_hd__o2111a_1 _8252_ (.A1(_3933_),
    .A2(_3398_),
    .B1(_3417_),
    .C1(_3447_),
    .D1(_3449_),
    .X(_3450_));
 sky130_fd_sc_hd__a31o_1 _8253_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3446_),
    .B1(_3450_),
    .X(net94));
 sky130_fd_sc_hd__nor2_1 _8254_ (.A(_3257_),
    .B(_3259_),
    .Y(_3451_));
 sky130_fd_sc_hd__xnor2_1 _8255_ (.A(_3260_),
    .B(_3451_),
    .Y(_3452_));
 sky130_fd_sc_hd__mux2_1 _8256_ (.A0(_3445_),
    .A1(_3452_),
    .S(_3320_),
    .X(_3453_));
 sky130_fd_sc_hd__or2_1 _8257_ (.A(_3939_),
    .B(_3398_),
    .X(_3454_));
 sky130_fd_sc_hd__or3_1 _8258_ (.A(_3932_),
    .B(_3936_),
    .C(_3399_),
    .X(_3455_));
 sky130_fd_sc_hd__o2111a_1 _8259_ (.A1(_3933_),
    .A2(_3395_),
    .B1(_3417_),
    .C1(_3454_),
    .D1(_3455_),
    .X(_3456_));
 sky130_fd_sc_hd__a31o_1 _8260_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3453_),
    .B1(_3456_),
    .X(net95));
 sky130_fd_sc_hd__and2_1 _8261_ (.A(_3262_),
    .B(_3263_),
    .X(_3458_));
 sky130_fd_sc_hd__xnor2_2 _8262_ (.A(_3264_),
    .B(_3458_),
    .Y(_3459_));
 sky130_fd_sc_hd__mux2_1 _8263_ (.A0(_3452_),
    .A1(_3459_),
    .S(_3320_),
    .X(_3460_));
 sky130_fd_sc_hd__or3_1 _8264_ (.A(_3932_),
    .B(_3936_),
    .C(_3398_),
    .X(_3461_));
 sky130_fd_sc_hd__o21a_1 _8265_ (.A1(_3933_),
    .A2(_3394_),
    .B1(_3461_),
    .X(_3462_));
 sky130_fd_sc_hd__o211a_1 _8266_ (.A1(_3939_),
    .A2(_3395_),
    .B1(_3417_),
    .C1(_3462_),
    .X(_3463_));
 sky130_fd_sc_hd__a31o_1 _8267_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3460_),
    .B1(_3463_),
    .X(net96));
 sky130_fd_sc_hd__nand2_1 _8268_ (.A(_3266_),
    .B(_3268_),
    .Y(_3464_));
 sky130_fd_sc_hd__xnor2_1 _8269_ (.A(_3269_),
    .B(_3464_),
    .Y(_3465_));
 sky130_fd_sc_hd__mux2_1 _8270_ (.A0(_3459_),
    .A1(_3465_),
    .S(_3320_),
    .X(_3466_));
 sky130_fd_sc_hd__or2_1 _8271_ (.A(_3939_),
    .B(_3394_),
    .X(_3468_));
 sky130_fd_sc_hd__or3_1 _8272_ (.A(_3932_),
    .B(_3936_),
    .C(_3395_),
    .X(_3469_));
 sky130_fd_sc_hd__o2111a_1 _8273_ (.A1(_3933_),
    .A2(_3392_),
    .B1(_3417_),
    .C1(_3468_),
    .D1(_3469_),
    .X(_3470_));
 sky130_fd_sc_hd__a31o_1 _8274_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3466_),
    .B1(_3470_),
    .X(net97));
 sky130_fd_sc_hd__and2_1 _8275_ (.A(_3271_),
    .B(_3272_),
    .X(_3471_));
 sky130_fd_sc_hd__xnor2_1 _8276_ (.A(_3273_),
    .B(_3471_),
    .Y(_3472_));
 sky130_fd_sc_hd__mux2_1 _8277_ (.A0(_3465_),
    .A1(_3472_),
    .S(_3320_),
    .X(_3473_));
 sky130_fd_sc_hd__or2_1 _8278_ (.A(_3939_),
    .B(_3392_),
    .X(_3474_));
 sky130_fd_sc_hd__nand2_1 _8279_ (.A(_3932_),
    .B(_3391_),
    .Y(_3475_));
 sky130_fd_sc_hd__o311a_1 _8280_ (.A1(_3932_),
    .A2(_3936_),
    .A3(_3394_),
    .B1(_3417_),
    .C1(_3475_),
    .X(_3476_));
 sky130_fd_sc_hd__a32o_1 _8281_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3473_),
    .B1(_3474_),
    .B2(_3476_),
    .X(net67));
 sky130_fd_sc_hd__nand2_1 _8282_ (.A(_3275_),
    .B(_3276_),
    .Y(_3478_));
 sky130_fd_sc_hd__xnor2_1 _8283_ (.A(_3277_),
    .B(_3478_),
    .Y(_3479_));
 sky130_fd_sc_hd__mux2_1 _8284_ (.A0(_3472_),
    .A1(_3479_),
    .S(_3320_),
    .X(_3480_));
 sky130_fd_sc_hd__nand2_1 _8285_ (.A(_3938_),
    .B(_3391_),
    .Y(_3481_));
 sky130_fd_sc_hd__nand2_1 _8286_ (.A(_3932_),
    .B(_3389_),
    .Y(_3482_));
 sky130_fd_sc_hd__o311a_1 _8287_ (.A1(_3932_),
    .A2(_3936_),
    .A3(_3392_),
    .B1(_3417_),
    .C1(_3482_),
    .X(_3483_));
 sky130_fd_sc_hd__a32o_1 _8288_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3480_),
    .B1(_3481_),
    .B2(_3483_),
    .X(net68));
 sky130_fd_sc_hd__and2_1 _8289_ (.A(_3280_),
    .B(_3281_),
    .X(_3484_));
 sky130_fd_sc_hd__xnor2_1 _8290_ (.A(_3282_),
    .B(_3484_),
    .Y(_3485_));
 sky130_fd_sc_hd__mux2_1 _8291_ (.A0(_3479_),
    .A1(_3485_),
    .S(_3320_),
    .X(_3487_));
 sky130_fd_sc_hd__mux2_1 _8292_ (.A0(_3389_),
    .A1(_3391_),
    .S(_3937_),
    .X(_3488_));
 sky130_fd_sc_hd__mux2_1 _8293_ (.A0(_3488_),
    .A1(_3388_),
    .S(_3932_),
    .X(_3489_));
 sky130_fd_sc_hd__inv_2 _8294_ (.A(_3489_),
    .Y(_3490_));
 sky130_fd_sc_hd__a32o_1 _8295_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3487_),
    .B1(_3490_),
    .B2(_3417_),
    .X(net69));
 sky130_fd_sc_hd__nand2_1 _8296_ (.A(_3284_),
    .B(_3285_),
    .Y(_3491_));
 sky130_fd_sc_hd__xor2_1 _8297_ (.A(_3286_),
    .B(_3491_),
    .X(_3492_));
 sky130_fd_sc_hd__mux2_1 _8298_ (.A0(_3485_),
    .A1(_3492_),
    .S(_3320_),
    .X(_3493_));
 sky130_fd_sc_hd__mux2_1 _8299_ (.A0(_3388_),
    .A1(_3389_),
    .S(_3937_),
    .X(_3494_));
 sky130_fd_sc_hd__mux2_1 _8300_ (.A0(_3494_),
    .A1(_3385_),
    .S(_3932_),
    .X(_3495_));
 sky130_fd_sc_hd__inv_2 _8301_ (.A(_3495_),
    .Y(_3497_));
 sky130_fd_sc_hd__a32o_1 _8302_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3493_),
    .B1(_3497_),
    .B2(_3417_),
    .X(net70));
 sky130_fd_sc_hd__and2_1 _8303_ (.A(_3288_),
    .B(_3290_),
    .X(_3498_));
 sky130_fd_sc_hd__xnor2_1 _8304_ (.A(_3291_),
    .B(_3498_),
    .Y(_3499_));
 sky130_fd_sc_hd__mux2_1 _8305_ (.A0(_3492_),
    .A1(_3499_),
    .S(_3320_),
    .X(_3500_));
 sky130_fd_sc_hd__and3_1 _8306_ (.A(_3933_),
    .B(_3937_),
    .C(_3388_),
    .X(_3501_));
 sky130_fd_sc_hd__a221oi_1 _8307_ (.A1(_3932_),
    .A2(_3383_),
    .B1(_3385_),
    .B2(_3938_),
    .C1(_3501_),
    .Y(_3502_));
 sky130_fd_sc_hd__a32o_1 _8308_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3500_),
    .B1(_3502_),
    .B2(_3417_),
    .X(net71));
 sky130_fd_sc_hd__nand2_1 _8309_ (.A(_3184_),
    .B(_3185_),
    .Y(_3503_));
 sky130_fd_sc_hd__xnor2_1 _8310_ (.A(_3293_),
    .B(_3503_),
    .Y(_3504_));
 sky130_fd_sc_hd__mux2_1 _8311_ (.A0(_3499_),
    .A1(_3504_),
    .S(_3320_),
    .X(_3506_));
 sky130_fd_sc_hd__mux2_1 _8312_ (.A0(_3383_),
    .A1(_3385_),
    .S(_3937_),
    .X(_3507_));
 sky130_fd_sc_hd__mux2_1 _8313_ (.A0(_3507_),
    .A1(_3381_),
    .S(_3932_),
    .X(_3508_));
 sky130_fd_sc_hd__inv_2 _8314_ (.A(_3508_),
    .Y(_3509_));
 sky130_fd_sc_hd__a32o_1 _8315_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3506_),
    .B1(_3509_),
    .B2(_3417_),
    .X(net72));
 sky130_fd_sc_hd__nand2_1 _8316_ (.A(_3295_),
    .B(_3296_),
    .Y(_3510_));
 sky130_fd_sc_hd__xnor2_1 _8317_ (.A(_3298_),
    .B(_3510_),
    .Y(_3511_));
 sky130_fd_sc_hd__mux2_1 _8318_ (.A0(_3504_),
    .A1(_3511_),
    .S(_3320_),
    .X(_3512_));
 sky130_fd_sc_hd__mux2_1 _8319_ (.A0(_3381_),
    .A1(_3383_),
    .S(_3937_),
    .X(_3513_));
 sky130_fd_sc_hd__mux2_1 _8320_ (.A0(_3513_),
    .A1(_3379_),
    .S(_3932_),
    .X(_3514_));
 sky130_fd_sc_hd__inv_2 _8321_ (.A(_3514_),
    .Y(_3516_));
 sky130_fd_sc_hd__a32o_1 _8322_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3512_),
    .B1(_3516_),
    .B2(_3417_),
    .X(net73));
 sky130_fd_sc_hd__and2_1 _8323_ (.A(_3176_),
    .B(_3177_),
    .X(_3517_));
 sky130_fd_sc_hd__xor2_1 _8324_ (.A(_3301_),
    .B(_3517_),
    .X(_3518_));
 sky130_fd_sc_hd__inv_2 _8325_ (.A(_3518_),
    .Y(_3519_));
 sky130_fd_sc_hd__mux2_1 _8326_ (.A0(_3511_),
    .A1(_3519_),
    .S(_3320_),
    .X(_3520_));
 sky130_fd_sc_hd__mux2_1 _8327_ (.A0(_3379_),
    .A1(_3381_),
    .S(_3937_),
    .X(_3521_));
 sky130_fd_sc_hd__mux2_1 _8328_ (.A0(_3521_),
    .A1(_3377_),
    .S(_3932_),
    .X(_3522_));
 sky130_fd_sc_hd__inv_2 _8329_ (.A(_3522_),
    .Y(_3523_));
 sky130_fd_sc_hd__a32o_1 _8330_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3520_),
    .B1(_3523_),
    .B2(_3417_),
    .X(net74));
 sky130_fd_sc_hd__nand2_1 _8331_ (.A(_3303_),
    .B(_3304_),
    .Y(_3525_));
 sky130_fd_sc_hd__xnor2_1 _8332_ (.A(_3305_),
    .B(_3525_),
    .Y(_3526_));
 sky130_fd_sc_hd__mux2_1 _8333_ (.A0(_3518_),
    .A1(_3526_),
    .S(_3320_),
    .X(_3527_));
 sky130_fd_sc_hd__inv_2 _8334_ (.A(_3527_),
    .Y(_3528_));
 sky130_fd_sc_hd__mux2_1 _8335_ (.A0(_3377_),
    .A1(_3379_),
    .S(_3937_),
    .X(_3529_));
 sky130_fd_sc_hd__mux2_1 _8336_ (.A0(_3529_),
    .A1(_3374_),
    .S(_3932_),
    .X(_3530_));
 sky130_fd_sc_hd__inv_2 _8337_ (.A(_3530_),
    .Y(_3531_));
 sky130_fd_sc_hd__a32o_1 _8338_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3528_),
    .B1(_3531_),
    .B2(_3417_),
    .X(net75));
 sky130_fd_sc_hd__and2_1 _8339_ (.A(_3170_),
    .B(_3171_),
    .X(_3532_));
 sky130_fd_sc_hd__xor2_1 _8340_ (.A(_3307_),
    .B(_3532_),
    .X(_3533_));
 sky130_fd_sc_hd__inv_2 _8341_ (.A(_3533_),
    .Y(_3535_));
 sky130_fd_sc_hd__mux2_1 _8342_ (.A0(_3526_),
    .A1(_3533_),
    .S(_3320_),
    .X(_3536_));
 sky130_fd_sc_hd__inv_2 _8343_ (.A(_3536_),
    .Y(_3537_));
 sky130_fd_sc_hd__and3_1 _8344_ (.A(_3933_),
    .B(_3937_),
    .C(_3377_),
    .X(_3538_));
 sky130_fd_sc_hd__a221oi_1 _8345_ (.A1(_3932_),
    .A2(_3373_),
    .B1(_3374_),
    .B2(_3938_),
    .C1(_3538_),
    .Y(_3539_));
 sky130_fd_sc_hd__a32o_1 _8346_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3537_),
    .B1(_3539_),
    .B2(_3417_),
    .X(net76));
 sky130_fd_sc_hd__nand2_1 _8347_ (.A(_3312_),
    .B(_3313_),
    .Y(_3540_));
 sky130_fd_sc_hd__xnor2_1 _8348_ (.A(_3315_),
    .B(_3540_),
    .Y(_3541_));
 sky130_fd_sc_hd__mux2_1 _8349_ (.A0(_3535_),
    .A1(_3541_),
    .S(_3320_),
    .X(_3542_));
 sky130_fd_sc_hd__mux2_1 _8350_ (.A0(_3373_),
    .A1(_3374_),
    .S(_3937_),
    .X(_3543_));
 sky130_fd_sc_hd__mux2_1 _8351_ (.A0(_3543_),
    .A1(_3371_),
    .S(_3932_),
    .X(_3545_));
 sky130_fd_sc_hd__inv_2 _8352_ (.A(_3545_),
    .Y(_3546_));
 sky130_fd_sc_hd__a32o_1 _8353_ (.A1(_3346_),
    .A2(_3351_),
    .A3(_3542_),
    .B1(_3546_),
    .B2(_3417_),
    .X(net78));
 sky130_fd_sc_hd__nand2_1 _8354_ (.A(_3165_),
    .B(_3166_),
    .Y(_3547_));
 sky130_fd_sc_hd__xor2_1 _8355_ (.A(_3317_),
    .B(_3547_),
    .X(_3548_));
 sky130_fd_sc_hd__or2_1 _8356_ (.A(_3320_),
    .B(_3541_),
    .X(_3549_));
 sky130_fd_sc_hd__a21oi_1 _8357_ (.A1(_3320_),
    .A2(_3548_),
    .B1(_3350_),
    .Y(_3550_));
 sky130_fd_sc_hd__and3_1 _8358_ (.A(_3933_),
    .B(_3937_),
    .C(_3373_),
    .X(_3551_));
 sky130_fd_sc_hd__a221oi_1 _8359_ (.A1(_3938_),
    .A2(_3371_),
    .B1(_3415_),
    .B2(_3932_),
    .C1(_3551_),
    .Y(_3552_));
 sky130_fd_sc_hd__a32o_1 _8360_ (.A1(_3346_),
    .A2(_3549_),
    .A3(_3550_),
    .B1(_3552_),
    .B2(_3417_),
    .X(net79));
 sky130_fd_sc_hd__o22a_1 _8361_ (.A1(_3161_),
    .A2(_3319_),
    .B1(_3320_),
    .B2(_3548_),
    .X(_3554_));
 sky130_fd_sc_hd__nor2_1 _8362_ (.A(_3350_),
    .B(_3554_),
    .Y(_3555_));
 sky130_fd_sc_hd__a31o_1 _8363_ (.A1(_3342_),
    .A2(_3345_),
    .A3(_3555_),
    .B1(_3946_),
    .X(_3556_));
 sky130_fd_sc_hd__o21ai_1 _8364_ (.A1(_3932_),
    .A2(_3371_),
    .B1(_3937_),
    .Y(_3557_));
 sky130_fd_sc_hd__nand2_1 _8365_ (.A(_3938_),
    .B(_3415_),
    .Y(_3558_));
 sky130_fd_sc_hd__a32o_1 _8366_ (.A1(_3417_),
    .A2(_3557_),
    .A3(_3558_),
    .B1(_3556_),
    .B2(net65),
    .X(net80));
 sky130_fd_sc_hd__nand2_1 _8367_ (.A(_3335_),
    .B(_3351_),
    .Y(_3559_));
 sky130_fd_sc_hd__a21o_1 _8368_ (.A1(_3342_),
    .A2(_3559_),
    .B1(_3343_),
    .X(_3560_));
 sky130_fd_sc_hd__and3_4 _8369_ (.A(_0308_),
    .B(_0451_),
    .C(_3947_),
    .X(_3561_));
 sky130_fd_sc_hd__mux2_1 _8370_ (.A0(net16),
    .A1(net48),
    .S(_0858_),
    .X(_3562_));
 sky130_fd_sc_hd__nor2_1 _8371_ (.A(_3939_),
    .B(_3562_),
    .Y(_3564_));
 sky130_fd_sc_hd__a211o_1 _8372_ (.A1(_3939_),
    .A2(_3562_),
    .B1(_3564_),
    .C1(_3416_),
    .X(_3565_));
 sky130_fd_sc_hd__a22oi_2 _8373_ (.A1(_3560_),
    .A2(_3561_),
    .B1(_3565_),
    .B2(_1122_),
    .Y(net81));
 sky130_fd_sc_hd__mux2_1 _8374_ (.A0(net17),
    .A1(net49),
    .S(_0858_),
    .X(_3566_));
 sky130_fd_sc_hd__nand2_1 _8375_ (.A(_3936_),
    .B(_3566_),
    .Y(_3567_));
 sky130_fd_sc_hd__nand2_1 _8376_ (.A(_3562_),
    .B(_3566_),
    .Y(_3568_));
 sky130_fd_sc_hd__or2_1 _8377_ (.A(_3562_),
    .B(_3566_),
    .X(_3569_));
 sky130_fd_sc_hd__nand2_1 _8378_ (.A(_3568_),
    .B(_3569_),
    .Y(_3570_));
 sky130_fd_sc_hd__a21oi_1 _8379_ (.A1(_3937_),
    .A2(_3570_),
    .B1(_3932_),
    .Y(_3571_));
 sky130_fd_sc_hd__a22o_1 _8380_ (.A1(_3932_),
    .A2(_3570_),
    .B1(_3571_),
    .B2(_3567_),
    .X(_3572_));
 sky130_fd_sc_hd__o21a_1 _8381_ (.A1(_3416_),
    .A2(_3572_),
    .B1(_1122_),
    .X(_3574_));
 sky130_fd_sc_hd__a21oi_1 _8382_ (.A1(_0638_),
    .A2(_3320_),
    .B1(_3972_),
    .Y(_3575_));
 sky130_fd_sc_hd__a211o_1 _8383_ (.A1(_3320_),
    .A2(_3321_),
    .B1(_3350_),
    .C1(_3575_),
    .X(_3576_));
 sky130_fd_sc_hd__a21o_1 _8384_ (.A1(_3342_),
    .A2(_3576_),
    .B1(_3343_),
    .X(_3577_));
 sky130_fd_sc_hd__a21oi_1 _8385_ (.A1(_3561_),
    .A2(_3577_),
    .B1(_3574_),
    .Y(net82));
 sky130_fd_sc_hd__mux2_1 _8386_ (.A0(net18),
    .A1(net50),
    .S(_0858_),
    .X(_3578_));
 sky130_fd_sc_hd__or2_1 _8387_ (.A(_3936_),
    .B(_3569_),
    .X(_3579_));
 sky130_fd_sc_hd__mux2_1 _8388_ (.A0(_3579_),
    .A1(_3568_),
    .S(_3932_),
    .X(_3580_));
 sky130_fd_sc_hd__xor2_1 _8389_ (.A(_3578_),
    .B(_3580_),
    .X(_3581_));
 sky130_fd_sc_hd__o21a_1 _8390_ (.A1(_3416_),
    .A2(_3581_),
    .B1(_1122_),
    .X(_3582_));
 sky130_fd_sc_hd__a21oi_1 _8391_ (.A1(_3320_),
    .A2(_3321_),
    .B1(_3323_),
    .Y(_3584_));
 sky130_fd_sc_hd__a31o_1 _8392_ (.A1(_3320_),
    .A2(_3321_),
    .A3(_3323_),
    .B1(_3350_),
    .X(_3585_));
 sky130_fd_sc_hd__or2_1 _8393_ (.A(_3584_),
    .B(_3585_),
    .X(_3586_));
 sky130_fd_sc_hd__a21o_1 _8394_ (.A1(_3342_),
    .A2(_3586_),
    .B1(_3343_),
    .X(_3587_));
 sky130_fd_sc_hd__a21oi_1 _8395_ (.A1(_3561_),
    .A2(_3587_),
    .B1(_3582_),
    .Y(net83));
 sky130_fd_sc_hd__nand3b_1 _8396_ (.A_N(_3325_),
    .B(_3340_),
    .C(_3351_),
    .Y(_3588_));
 sky130_fd_sc_hd__a21o_1 _8397_ (.A1(_3342_),
    .A2(_3588_),
    .B1(_3343_),
    .X(_3589_));
 sky130_fd_sc_hd__mux2_2 _8398_ (.A0(net19),
    .A1(net51),
    .S(_0858_),
    .X(_3590_));
 sky130_fd_sc_hd__and3_1 _8399_ (.A(_3562_),
    .B(_3566_),
    .C(_3578_),
    .X(_3591_));
 sky130_fd_sc_hd__or2_1 _8400_ (.A(_3578_),
    .B(_3579_),
    .X(_3592_));
 sky130_fd_sc_hd__inv_2 _8401_ (.A(_3592_),
    .Y(_3594_));
 sky130_fd_sc_hd__mux2_1 _8402_ (.A0(_3591_),
    .A1(_3594_),
    .S(_3933_),
    .X(_3595_));
 sky130_fd_sc_hd__a21oi_1 _8403_ (.A1(_3590_),
    .A2(_3595_),
    .B1(_3416_),
    .Y(_3596_));
 sky130_fd_sc_hd__and2_1 _8404_ (.A(_3590_),
    .B(_3591_),
    .X(_3597_));
 sky130_fd_sc_hd__nor2_1 _8405_ (.A(_3590_),
    .B(_3592_),
    .Y(_3598_));
 sky130_fd_sc_hd__o21ai_1 _8406_ (.A1(_3590_),
    .A2(_3595_),
    .B1(_3596_),
    .Y(_3599_));
 sky130_fd_sc_hd__a22oi_2 _8407_ (.A1(_3561_),
    .A2(_3589_),
    .B1(_3599_),
    .B2(_1122_),
    .Y(net84));
 sky130_fd_sc_hd__mux2_2 _8408_ (.A0(net20),
    .A1(net52),
    .S(_0803_),
    .X(_3600_));
 sky130_fd_sc_hd__mux2_1 _8409_ (.A0(_3597_),
    .A1(_3598_),
    .S(_3933_),
    .X(_3601_));
 sky130_fd_sc_hd__a21oi_1 _8410_ (.A1(_3600_),
    .A2(_3601_),
    .B1(_3416_),
    .Y(_3602_));
 sky130_fd_sc_hd__o21ai_1 _8411_ (.A1(_3600_),
    .A2(_3601_),
    .B1(_3602_),
    .Y(_3604_));
 sky130_fd_sc_hd__a21oi_1 _8412_ (.A1(_3325_),
    .A2(_3330_),
    .B1(_3350_),
    .Y(_3605_));
 sky130_fd_sc_hd__o21ai_1 _8413_ (.A1(_3325_),
    .A2(_3330_),
    .B1(_3605_),
    .Y(_3606_));
 sky130_fd_sc_hd__a21o_1 _8414_ (.A1(_3342_),
    .A2(_3606_),
    .B1(_3343_),
    .X(_3607_));
 sky130_fd_sc_hd__a22oi_2 _8415_ (.A1(_1122_),
    .A2(_3604_),
    .B1(_3607_),
    .B2(_3561_),
    .Y(net85));
 sky130_fd_sc_hd__and3_1 _8416_ (.A(_3325_),
    .B(_3330_),
    .C(_3332_),
    .X(_3608_));
 sky130_fd_sc_hd__o21ai_1 _8417_ (.A1(_3334_),
    .A2(_3608_),
    .B1(_3351_),
    .Y(_3609_));
 sky130_fd_sc_hd__a21o_1 _8418_ (.A1(_3342_),
    .A2(_3609_),
    .B1(_3343_),
    .X(_3610_));
 sky130_fd_sc_hd__mux2_1 _8419_ (.A0(net21),
    .A1(net53),
    .S(_0858_),
    .X(_3611_));
 sky130_fd_sc_hd__o31ai_1 _8420_ (.A1(_3590_),
    .A2(_3592_),
    .A3(_3600_),
    .B1(_3611_),
    .Y(_3612_));
 sky130_fd_sc_hd__o41a_1 _8421_ (.A1(_3590_),
    .A2(_3592_),
    .A3(_3600_),
    .A4(_3611_),
    .B1(_3933_),
    .X(_3614_));
 sky130_fd_sc_hd__nand3_1 _8422_ (.A(_3597_),
    .B(_3600_),
    .C(_3611_),
    .Y(_3615_));
 sky130_fd_sc_hd__a31o_1 _8423_ (.A1(_3590_),
    .A2(_3591_),
    .A3(_3600_),
    .B1(_3611_),
    .X(_3616_));
 sky130_fd_sc_hd__nand2_1 _8424_ (.A(_3615_),
    .B(_3616_),
    .Y(_3617_));
 sky130_fd_sc_hd__a22o_1 _8425_ (.A1(_3612_),
    .A2(_3614_),
    .B1(_3617_),
    .B2(_3932_),
    .X(_3618_));
 sky130_fd_sc_hd__o21a_1 _8426_ (.A1(_3416_),
    .A2(_3618_),
    .B1(_1122_),
    .X(_3619_));
 sky130_fd_sc_hd__a21oi_1 _8427_ (.A1(_3561_),
    .A2(_3610_),
    .B1(_3619_),
    .Y(net86));
 sky130_fd_sc_hd__a21oi_2 _8428_ (.A1(_3932_),
    .A2(_3615_),
    .B1(_3614_),
    .Y(_3620_));
 sky130_fd_sc_hd__mux2_1 _8429_ (.A0(net22),
    .A1(net54),
    .S(_0803_),
    .X(_3621_));
 sky130_fd_sc_hd__nor2_1 _8430_ (.A(_3620_),
    .B(_3621_),
    .Y(_3622_));
 sky130_fd_sc_hd__a21o_1 _8431_ (.A1(_3620_),
    .A2(_3621_),
    .B1(_3416_),
    .X(_3624_));
 sky130_fd_sc_hd__o21a_1 _8432_ (.A1(_3622_),
    .A2(_3624_),
    .B1(_1122_),
    .X(_3625_));
 sky130_fd_sc_hd__or3_1 _8433_ (.A(_3327_),
    .B(_3328_),
    .C(_3350_),
    .X(_3626_));
 sky130_fd_sc_hd__a21o_1 _8434_ (.A1(_3342_),
    .A2(_3626_),
    .B1(_3343_),
    .X(_3627_));
 sky130_fd_sc_hd__a21oi_1 _8435_ (.A1(_3561_),
    .A2(_3627_),
    .B1(_3625_),
    .Y(net87));
 sky130_fd_sc_hd__xnor2_1 _8436_ (.A(_3932_),
    .B(_3621_),
    .Y(_3628_));
 sky130_fd_sc_hd__a21oi_1 _8437_ (.A1(_3620_),
    .A2(_3628_),
    .B1(_3349_),
    .Y(_3629_));
 sky130_fd_sc_hd__a311o_1 _8438_ (.A1(_3349_),
    .A2(_3620_),
    .A3(_3628_),
    .B1(_3629_),
    .C1(_3416_),
    .X(_3630_));
 sky130_fd_sc_hd__and4_1 _8439_ (.A(_3970_),
    .B(_3325_),
    .C(_3326_),
    .D(_3337_),
    .X(_3631_));
 sky130_fd_sc_hd__a31o_1 _8440_ (.A1(_3970_),
    .A2(_3325_),
    .A3(_3326_),
    .B1(_3337_),
    .X(_3632_));
 sky130_fd_sc_hd__or3b_1 _8441_ (.A(_3350_),
    .B(_3631_),
    .C_N(_3632_),
    .X(_3634_));
 sky130_fd_sc_hd__a21o_1 _8442_ (.A1(_3342_),
    .A2(_3634_),
    .B1(_3343_),
    .X(_3635_));
 sky130_fd_sc_hd__a22oi_2 _8443_ (.A1(_1122_),
    .A2(_3630_),
    .B1(_3635_),
    .B2(_3561_),
    .Y(net89));
 sky130_fd_sc_hd__mux2_1 _8444_ (.A0(net25),
    .A1(net57),
    .S(_3744_),
    .X(_3636_));
 sky130_fd_sc_hd__and2b_1 _8445_ (.A_N(_3416_),
    .B(_3636_),
    .X(_3637_));
 sky130_fd_sc_hd__mux2_1 _8446_ (.A0(net25),
    .A1(net57),
    .S(_0451_),
    .X(_3638_));
 sky130_fd_sc_hd__and4_1 _8447_ (.A(_0176_),
    .B(_1111_),
    .C(_3941_),
    .D(_3638_),
    .X(_3639_));
 sky130_fd_sc_hd__o22a_1 _8448_ (.A1(_0462_),
    .A2(_3637_),
    .B1(_3639_),
    .B2(_1122_),
    .X(_3640_));
 sky130_fd_sc_hd__a41o_1 _8449_ (.A1(_3745_),
    .A2(_3944_),
    .A3(_3945_),
    .A4(_3947_),
    .B1(_3640_),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_16 input1 (.A(in1[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_12 input2 (.A(in1[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_12 input3 (.A(in1[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_12 input4 (.A(in1[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_12 input5 (.A(in1[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_12 input6 (.A(in1[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_12 input7 (.A(in1[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_16 input8 (.A(in1[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_12 input9 (.A(in1[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 input10 (.A(in1[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_16 input11 (.A(in1[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_12 input12 (.A(in1[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_16 input13 (.A(in1[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_16 input14 (.A(in1[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_16 input15 (.A(in1[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(in1[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(in1[24]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(in1[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(in1[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in1[27]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(in1[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in1[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_12 input23 (.A(in1[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(in1[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(in1[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_12 input26 (.A(in1[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_12 input27 (.A(in1[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_12 input28 (.A(in1[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_12 input29 (.A(in1[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_12 input30 (.A(in1[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_12 input31 (.A(in1[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_16 input32 (.A(in1[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_12 input33 (.A(in2[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_16 input34 (.A(in2[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_8 input35 (.A(in2[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_12 input36 (.A(in2[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_12 input37 (.A(in2[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_8 input38 (.A(in2[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_16 input39 (.A(in2[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_8 input40 (.A(in2[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_8 input41 (.A(in2[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_8 input42 (.A(in2[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_12 input43 (.A(in2[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_12 input44 (.A(in2[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_16 input45 (.A(in2[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_16 input46 (.A(in2[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_16 input47 (.A(in2[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(in2[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(in2[24]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(in2[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(in2[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(in2[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(in2[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in2[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_12 input55 (.A(in2[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(in2[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(in2[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_12 input58 (.A(in2[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_12 input59 (.A(in2[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_12 input60 (.A(in2[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_12 input61 (.A(in2[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_12 input62 (.A(in2[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_16 input63 (.A(in2[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_12 input64 (.A(in2[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(sel),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_16 output66 (.A(net66),
    .X(result[0]));
 sky130_fd_sc_hd__clkbuf_16 output67 (.A(net67),
    .X(result[10]));
 sky130_fd_sc_hd__clkbuf_16 output68 (.A(net68),
    .X(result[11]));
 sky130_fd_sc_hd__clkbuf_16 output69 (.A(net69),
    .X(result[12]));
 sky130_fd_sc_hd__clkbuf_16 output70 (.A(net70),
    .X(result[13]));
 sky130_fd_sc_hd__clkbuf_16 output71 (.A(net71),
    .X(result[14]));
 sky130_fd_sc_hd__clkbuf_16 output72 (.A(net72),
    .X(result[15]));
 sky130_fd_sc_hd__clkbuf_16 output73 (.A(net73),
    .X(result[16]));
 sky130_fd_sc_hd__clkbuf_16 output74 (.A(net74),
    .X(result[17]));
 sky130_fd_sc_hd__clkbuf_16 output75 (.A(net75),
    .X(result[18]));
 sky130_fd_sc_hd__clkbuf_16 output76 (.A(net76),
    .X(result[19]));
 sky130_fd_sc_hd__clkbuf_16 output77 (.A(net77),
    .X(result[1]));
 sky130_fd_sc_hd__clkbuf_16 output78 (.A(net78),
    .X(result[20]));
 sky130_fd_sc_hd__clkbuf_16 output79 (.A(net79),
    .X(result[21]));
 sky130_fd_sc_hd__clkbuf_16 output80 (.A(net80),
    .X(result[22]));
 sky130_fd_sc_hd__clkbuf_16 output81 (.A(net81),
    .X(result[23]));
 sky130_fd_sc_hd__clkbuf_16 output82 (.A(net82),
    .X(result[24]));
 sky130_fd_sc_hd__clkbuf_16 output83 (.A(net83),
    .X(result[25]));
 sky130_fd_sc_hd__clkbuf_16 output84 (.A(net84),
    .X(result[26]));
 sky130_fd_sc_hd__clkbuf_16 output85 (.A(net85),
    .X(result[27]));
 sky130_fd_sc_hd__clkbuf_16 output86 (.A(net86),
    .X(result[28]));
 sky130_fd_sc_hd__clkbuf_16 output87 (.A(net87),
    .X(result[29]));
 sky130_fd_sc_hd__clkbuf_16 output88 (.A(net88),
    .X(result[2]));
 sky130_fd_sc_hd__clkbuf_16 output89 (.A(net89),
    .X(result[30]));
 sky130_fd_sc_hd__clkbuf_16 output90 (.A(net90),
    .X(result[31]));
 sky130_fd_sc_hd__clkbuf_16 output91 (.A(net91),
    .X(result[3]));
 sky130_fd_sc_hd__clkbuf_16 output92 (.A(net92),
    .X(result[4]));
 sky130_fd_sc_hd__clkbuf_16 output93 (.A(net93),
    .X(result[5]));
 sky130_fd_sc_hd__clkbuf_16 output94 (.A(net94),
    .X(result[6]));
 sky130_fd_sc_hd__clkbuf_16 output95 (.A(net95),
    .X(result[7]));
 sky130_fd_sc_hd__clkbuf_16 output96 (.A(net96),
    .X(result[8]));
 sky130_fd_sc_hd__clkbuf_16 output97 (.A(net97),
    .X(result[9]));
 sky130_fd_sc_hd__buf_8 max_cap98 (.A(_0814_),
    .X(net98));
endmodule
