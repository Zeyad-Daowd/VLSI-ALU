module booth_multiplier_route (clk,
    done,
    rst,
    start,
    M,
    Q,
    result);
 input clk;
 output done;
 input rst;
 input start;
 input [31:0] M;
 input [31:0] Q;
 output [63:0] result;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire \current_multiplier[0] ;
 wire \current_multiplier[10] ;
 wire \current_multiplier[11] ;
 wire \current_multiplier[12] ;
 wire \current_multiplier[13] ;
 wire \current_multiplier[14] ;
 wire \current_multiplier[15] ;
 wire \current_multiplier[16] ;
 wire \current_multiplier[17] ;
 wire \current_multiplier[18] ;
 wire \current_multiplier[19] ;
 wire \current_multiplier[1] ;
 wire \current_multiplier[20] ;
 wire \current_multiplier[21] ;
 wire \current_multiplier[22] ;
 wire \current_multiplier[23] ;
 wire \current_multiplier[24] ;
 wire \current_multiplier[25] ;
 wire \current_multiplier[26] ;
 wire \current_multiplier[27] ;
 wire \current_multiplier[28] ;
 wire \current_multiplier[29] ;
 wire \current_multiplier[2] ;
 wire \current_multiplier[30] ;
 wire \current_multiplier[31] ;
 wire \current_multiplier[3] ;
 wire \current_multiplier[4] ;
 wire \current_multiplier[5] ;
 wire \current_multiplier[6] ;
 wire \current_multiplier[7] ;
 wire \current_multiplier[8] ;
 wire \current_multiplier[9] ;
 wire \current_state[0] ;
 wire \current_state[1] ;
 wire \current_state[2] ;
 wire \extended_operand[0] ;
 wire \extended_operand[10] ;
 wire \extended_operand[11] ;
 wire \extended_operand[12] ;
 wire \extended_operand[13] ;
 wire \extended_operand[14] ;
 wire \extended_operand[15] ;
 wire \extended_operand[16] ;
 wire \extended_operand[17] ;
 wire \extended_operand[18] ;
 wire \extended_operand[19] ;
 wire \extended_operand[1] ;
 wire \extended_operand[20] ;
 wire \extended_operand[21] ;
 wire \extended_operand[22] ;
 wire \extended_operand[23] ;
 wire \extended_operand[24] ;
 wire \extended_operand[25] ;
 wire \extended_operand[26] ;
 wire \extended_operand[27] ;
 wire \extended_operand[28] ;
 wire \extended_operand[29] ;
 wire \extended_operand[2] ;
 wire \extended_operand[30] ;
 wire \extended_operand[31] ;
 wire \extended_operand[3] ;
 wire \extended_operand[4] ;
 wire \extended_operand[5] ;
 wire \extended_operand[6] ;
 wire \extended_operand[7] ;
 wire \extended_operand[8] ;
 wire \extended_operand[9] ;
 wire \iteration_count[0] ;
 wire \iteration_count[1] ;
 wire \iteration_count[2] ;
 wire \iteration_count[3] ;
 wire \iteration_count[4] ;
 wire \iteration_count[5] ;
 wire last_bit;
 wire \next_state[0] ;
 wire \next_state[1] ;
 wire \next_state[2] ;
 wire \partial_sum[0] ;
 wire \partial_sum[10] ;
 wire \partial_sum[11] ;
 wire \partial_sum[12] ;
 wire \partial_sum[13] ;
 wire \partial_sum[14] ;
 wire \partial_sum[15] ;
 wire \partial_sum[16] ;
 wire \partial_sum[17] ;
 wire \partial_sum[18] ;
 wire \partial_sum[19] ;
 wire \partial_sum[1] ;
 wire \partial_sum[20] ;
 wire \partial_sum[21] ;
 wire \partial_sum[22] ;
 wire \partial_sum[23] ;
 wire \partial_sum[24] ;
 wire \partial_sum[25] ;
 wire \partial_sum[26] ;
 wire \partial_sum[27] ;
 wire \partial_sum[28] ;
 wire \partial_sum[29] ;
 wire \partial_sum[2] ;
 wire \partial_sum[30] ;
 wire \partial_sum[31] ;
 wire \partial_sum[32] ;
 wire \partial_sum[33] ;
 wire \partial_sum[34] ;
 wire \partial_sum[35] ;
 wire \partial_sum[36] ;
 wire \partial_sum[37] ;
 wire \partial_sum[38] ;
 wire \partial_sum[39] ;
 wire \partial_sum[3] ;
 wire \partial_sum[40] ;
 wire \partial_sum[41] ;
 wire \partial_sum[42] ;
 wire \partial_sum[43] ;
 wire \partial_sum[44] ;
 wire \partial_sum[45] ;
 wire \partial_sum[46] ;
 wire \partial_sum[47] ;
 wire \partial_sum[48] ;
 wire \partial_sum[49] ;
 wire \partial_sum[4] ;
 wire \partial_sum[50] ;
 wire \partial_sum[51] ;
 wire \partial_sum[52] ;
 wire \partial_sum[53] ;
 wire \partial_sum[54] ;
 wire \partial_sum[55] ;
 wire \partial_sum[56] ;
 wire \partial_sum[57] ;
 wire \partial_sum[58] ;
 wire \partial_sum[59] ;
 wire \partial_sum[5] ;
 wire \partial_sum[60] ;
 wire \partial_sum[61] ;
 wire \partial_sum[62] ;
 wire \partial_sum[63] ;
 wire \partial_sum[6] ;
 wire \partial_sum[7] ;
 wire \partial_sum[8] ;
 wire \partial_sum[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__inv_2 _1056_ (.A(\current_multiplier[0] ),
    .Y(_0772_));
 sky130_fd_sc_hd__inv_2 _1057_ (.A(\partial_sum[27] ),
    .Y(_0773_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(\partial_sum[25] ),
    .Y(_0774_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(\partial_sum[23] ),
    .Y(_0775_));
 sky130_fd_sc_hd__inv_2 _1060_ (.A(\partial_sum[22] ),
    .Y(_0776_));
 sky130_fd_sc_hd__inv_2 _1061_ (.A(\partial_sum[18] ),
    .Y(_0777_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(\partial_sum[15] ),
    .Y(_0778_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(\partial_sum[10] ),
    .Y(_0779_));
 sky130_fd_sc_hd__inv_2 _1064_ (.A(\partial_sum[7] ),
    .Y(_0780_));
 sky130_fd_sc_hd__inv_2 _1065_ (.A(\partial_sum[6] ),
    .Y(_0781_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(\extended_operand[31] ),
    .Y(_0782_));
 sky130_fd_sc_hd__inv_2 _1067_ (.A(\extended_operand[18] ),
    .Y(_0783_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(net217),
    .Y(_0000_));
 sky130_fd_sc_hd__nor2_2 _1069_ (.A(\current_state[0] ),
    .B(\current_state[1] ),
    .Y(_0784_));
 sky130_fd_sc_hd__and2_1 _1070_ (.A(net212),
    .B(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__nand2_2 _1071_ (.A(\current_state[2] ),
    .B(_0784_),
    .Y(_0786_));
 sky130_fd_sc_hd__or3_1 _1072_ (.A(\iteration_count[2] ),
    .B(\iteration_count[1] ),
    .C(\iteration_count[0] ),
    .X(_0787_));
 sky130_fd_sc_hd__or2_1 _1073_ (.A(\iteration_count[3] ),
    .B(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__or3_1 _1074_ (.A(\iteration_count[5] ),
    .B(\iteration_count[4] ),
    .C(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__or4b_1 _1075_ (.A(\current_state[2] ),
    .B(\current_state[0] ),
    .C(\current_state[1] ),
    .D_N(net66),
    .X(_0790_));
 sky130_fd_sc_hd__o21ai_4 _1076_ (.A1(net212),
    .A2(net66),
    .B1(_0784_),
    .Y(_0791_));
 sky130_fd_sc_hd__o21a_1 _1077_ (.A1(\current_state[2] ),
    .A2(net66),
    .B1(_0784_),
    .X(_0792_));
 sky130_fd_sc_hd__o31ai_1 _1078_ (.A1(\iteration_count[4] ),
    .A2(_0788_),
    .A3(_0791_),
    .B1(\iteration_count[5] ),
    .Y(_0793_));
 sky130_fd_sc_hd__o211ai_1 _1079_ (.A1(net156),
    .A2(_0789_),
    .B1(net207),
    .C1(_0793_),
    .Y(_0402_));
 sky130_fd_sc_hd__xnor2_1 _1080_ (.A(\iteration_count[4] ),
    .B(_0788_),
    .Y(_0794_));
 sky130_fd_sc_hd__a22o_1 _1081_ (.A1(\iteration_count[4] ),
    .A2(_0791_),
    .B1(_0794_),
    .B2(net160),
    .X(_0401_));
 sky130_fd_sc_hd__nor2_1 _1082_ (.A(\iteration_count[0] ),
    .B(net156),
    .Y(_0795_));
 sky130_fd_sc_hd__nand2_1 _1083_ (.A(\iteration_count[3] ),
    .B(_0787_),
    .Y(_0796_));
 sky130_fd_sc_hd__nand2_1 _1084_ (.A(_0788_),
    .B(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__a22o_1 _1085_ (.A1(\iteration_count[3] ),
    .A2(_0791_),
    .B1(_0797_),
    .B2(net160),
    .X(_0400_));
 sky130_fd_sc_hd__o21ai_1 _1086_ (.A1(\iteration_count[1] ),
    .A2(\iteration_count[0] ),
    .B1(\iteration_count[2] ),
    .Y(_0798_));
 sky130_fd_sc_hd__nand2_1 _1087_ (.A(_0787_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__a22o_1 _1088_ (.A1(\iteration_count[2] ),
    .A2(_0791_),
    .B1(_0799_),
    .B2(net160),
    .X(_0399_));
 sky130_fd_sc_hd__a21o_1 _1089_ (.A1(\iteration_count[0] ),
    .A2(net212),
    .B1(_0791_),
    .X(_0800_));
 sky130_fd_sc_hd__mux2_1 _1090_ (.A0(_0795_),
    .A1(_0800_),
    .S(\iteration_count[1] ),
    .X(_0398_));
 sky130_fd_sc_hd__a21o_1 _1091_ (.A1(\iteration_count[0] ),
    .A2(_0791_),
    .B1(_0795_),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _1092_ (.A1(\current_multiplier[0] ),
    .A2(net160),
    .B1(_0791_),
    .B2(last_bit),
    .X(_0396_));
 sky130_fd_sc_hd__or2_1 _1093_ (.A(net57),
    .B(net203),
    .X(_0801_));
 sky130_fd_sc_hd__o221a_1 _1094_ (.A1(\partial_sum[0] ),
    .A2(net154),
    .B1(net150),
    .B2(\current_multiplier[31] ),
    .C1(_0801_),
    .X(_0395_));
 sky130_fd_sc_hd__or2_1 _1095_ (.A(net56),
    .B(net205),
    .X(_0802_));
 sky130_fd_sc_hd__o221a_1 _1096_ (.A1(\current_multiplier[31] ),
    .A2(net155),
    .B1(net151),
    .B2(\current_multiplier[30] ),
    .C1(_0802_),
    .X(_0394_));
 sky130_fd_sc_hd__or2_1 _1097_ (.A(net54),
    .B(net205),
    .X(_0803_));
 sky130_fd_sc_hd__o221a_1 _1098_ (.A1(\current_multiplier[30] ),
    .A2(net155),
    .B1(net151),
    .B2(\current_multiplier[29] ),
    .C1(_0803_),
    .X(_0393_));
 sky130_fd_sc_hd__or2_1 _1099_ (.A(net53),
    .B(net205),
    .X(_0804_));
 sky130_fd_sc_hd__o221a_1 _1100_ (.A1(\current_multiplier[29] ),
    .A2(net155),
    .B1(net151),
    .B2(\current_multiplier[28] ),
    .C1(_0804_),
    .X(_0392_));
 sky130_fd_sc_hd__or2_1 _1101_ (.A(net52),
    .B(net204),
    .X(_0805_));
 sky130_fd_sc_hd__o221a_1 _1102_ (.A1(\current_multiplier[28] ),
    .A2(net155),
    .B1(net151),
    .B2(\current_multiplier[27] ),
    .C1(_0805_),
    .X(_0391_));
 sky130_fd_sc_hd__or2_1 _1103_ (.A(net51),
    .B(net203),
    .X(_0806_));
 sky130_fd_sc_hd__o221a_1 _1104_ (.A1(\current_multiplier[27] ),
    .A2(net155),
    .B1(net151),
    .B2(\current_multiplier[26] ),
    .C1(_0806_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_1 _1105_ (.A(net50),
    .B(net202),
    .X(_0807_));
 sky130_fd_sc_hd__o221a_1 _1106_ (.A1(\current_multiplier[26] ),
    .A2(net154),
    .B1(net150),
    .B2(\current_multiplier[25] ),
    .C1(_0807_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_1 _1107_ (.A(net49),
    .B(net206),
    .X(_0808_));
 sky130_fd_sc_hd__o221a_1 _1108_ (.A1(\current_multiplier[25] ),
    .A2(net154),
    .B1(net150),
    .B2(\current_multiplier[24] ),
    .C1(_0808_),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _1109_ (.A(net48),
    .B(net202),
    .X(_0809_));
 sky130_fd_sc_hd__o221a_1 _1110_ (.A1(\current_multiplier[24] ),
    .A2(net154),
    .B1(net150),
    .B2(\current_multiplier[23] ),
    .C1(_0809_),
    .X(_0387_));
 sky130_fd_sc_hd__or2_1 _1111_ (.A(net47),
    .B(net202),
    .X(_0810_));
 sky130_fd_sc_hd__o221a_1 _1112_ (.A1(\current_multiplier[23] ),
    .A2(net154),
    .B1(net150),
    .B2(\current_multiplier[22] ),
    .C1(_0810_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _1113_ (.A(net46),
    .B(net202),
    .X(_0811_));
 sky130_fd_sc_hd__o221a_1 _1114_ (.A1(\current_multiplier[22] ),
    .A2(net154),
    .B1(net150),
    .B2(\current_multiplier[21] ),
    .C1(_0811_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _1115_ (.A(net45),
    .B(net203),
    .X(_0812_));
 sky130_fd_sc_hd__o221a_1 _1116_ (.A1(\current_multiplier[21] ),
    .A2(net154),
    .B1(net150),
    .B2(\current_multiplier[20] ),
    .C1(_0812_),
    .X(_0384_));
 sky130_fd_sc_hd__or2_1 _1117_ (.A(net43),
    .B(net203),
    .X(_0813_));
 sky130_fd_sc_hd__o221a_1 _1118_ (.A1(\current_multiplier[20] ),
    .A2(net154),
    .B1(net150),
    .B2(\current_multiplier[19] ),
    .C1(_0813_),
    .X(_0383_));
 sky130_fd_sc_hd__or2_1 _1119_ (.A(net42),
    .B(net203),
    .X(_0814_));
 sky130_fd_sc_hd__o221a_1 _1120_ (.A1(\current_multiplier[19] ),
    .A2(net154),
    .B1(net150),
    .B2(\current_multiplier[18] ),
    .C1(_0814_),
    .X(_0382_));
 sky130_fd_sc_hd__or2_1 _1121_ (.A(net41),
    .B(net202),
    .X(_0815_));
 sky130_fd_sc_hd__o221a_1 _1122_ (.A1(\current_multiplier[18] ),
    .A2(net154),
    .B1(net150),
    .B2(\current_multiplier[17] ),
    .C1(_0815_),
    .X(_0381_));
 sky130_fd_sc_hd__or2_1 _1123_ (.A(net40),
    .B(net204),
    .X(_0816_));
 sky130_fd_sc_hd__o221a_1 _1124_ (.A1(\current_multiplier[17] ),
    .A2(net155),
    .B1(net151),
    .B2(\current_multiplier[16] ),
    .C1(_0816_),
    .X(_0380_));
 sky130_fd_sc_hd__or2_1 _1125_ (.A(net39),
    .B(net204),
    .X(_0817_));
 sky130_fd_sc_hd__o221a_1 _1126_ (.A1(\current_multiplier[16] ),
    .A2(net155),
    .B1(net151),
    .B2(\current_multiplier[15] ),
    .C1(_0817_),
    .X(_0379_));
 sky130_fd_sc_hd__or2_1 _1127_ (.A(net38),
    .B(net204),
    .X(_0818_));
 sky130_fd_sc_hd__o221a_1 _1128_ (.A1(\current_multiplier[15] ),
    .A2(net156),
    .B1(net152),
    .B2(\current_multiplier[14] ),
    .C1(_0818_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_1 _1129_ (.A(net37),
    .B(net204),
    .X(_0819_));
 sky130_fd_sc_hd__o221a_1 _1130_ (.A1(\current_multiplier[14] ),
    .A2(net156),
    .B1(net152),
    .B2(\current_multiplier[13] ),
    .C1(_0819_),
    .X(_0377_));
 sky130_fd_sc_hd__or2_1 _1131_ (.A(net36),
    .B(net208),
    .X(_0820_));
 sky130_fd_sc_hd__o221a_1 _1132_ (.A1(\current_multiplier[13] ),
    .A2(net156),
    .B1(net152),
    .B2(\current_multiplier[12] ),
    .C1(_0820_),
    .X(_0376_));
 sky130_fd_sc_hd__or2_1 _1133_ (.A(net35),
    .B(net208),
    .X(_0821_));
 sky130_fd_sc_hd__o221a_1 _1134_ (.A1(\current_multiplier[12] ),
    .A2(net156),
    .B1(net152),
    .B2(\current_multiplier[11] ),
    .C1(_0821_),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _1135_ (.A(net34),
    .B(net208),
    .X(_0822_));
 sky130_fd_sc_hd__o221a_1 _1136_ (.A1(\current_multiplier[11] ),
    .A2(net157),
    .B1(net152),
    .B2(\current_multiplier[10] ),
    .C1(_0822_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_1 _1137_ (.A(net64),
    .B(net209),
    .X(_0823_));
 sky130_fd_sc_hd__o221a_1 _1138_ (.A1(\current_multiplier[10] ),
    .A2(net157),
    .B1(net152),
    .B2(\current_multiplier[9] ),
    .C1(_0823_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _1139_ (.A(net63),
    .B(net208),
    .X(_0824_));
 sky130_fd_sc_hd__o221a_1 _1140_ (.A1(\current_multiplier[9] ),
    .A2(net156),
    .B1(net152),
    .B2(\current_multiplier[8] ),
    .C1(_0824_),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _1141_ (.A(net62),
    .B(net210),
    .X(_0825_));
 sky130_fd_sc_hd__o221a_1 _1142_ (.A1(\current_multiplier[8] ),
    .A2(net156),
    .B1(net152),
    .B2(\current_multiplier[7] ),
    .C1(_0825_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _1143_ (.A(net61),
    .B(net210),
    .X(_0826_));
 sky130_fd_sc_hd__o221a_1 _1144_ (.A1(\current_multiplier[7] ),
    .A2(net157),
    .B1(net153),
    .B2(\current_multiplier[6] ),
    .C1(_0826_),
    .X(_0370_));
 sky130_fd_sc_hd__or2_1 _1145_ (.A(net60),
    .B(net209),
    .X(_0827_));
 sky130_fd_sc_hd__o221a_1 _1146_ (.A1(\current_multiplier[6] ),
    .A2(net157),
    .B1(net153),
    .B2(\current_multiplier[5] ),
    .C1(_0827_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_1 _1147_ (.A(net59),
    .B(net209),
    .X(_0828_));
 sky130_fd_sc_hd__o221a_1 _1148_ (.A1(\current_multiplier[5] ),
    .A2(net157),
    .B1(net153),
    .B2(\current_multiplier[4] ),
    .C1(_0828_),
    .X(_0368_));
 sky130_fd_sc_hd__or2_1 _1149_ (.A(net58),
    .B(net208),
    .X(_0829_));
 sky130_fd_sc_hd__o221a_1 _1150_ (.A1(\current_multiplier[4] ),
    .A2(net157),
    .B1(net153),
    .B2(\current_multiplier[3] ),
    .C1(_0829_),
    .X(_0367_));
 sky130_fd_sc_hd__or2_1 _1151_ (.A(net55),
    .B(net208),
    .X(_0830_));
 sky130_fd_sc_hd__o221a_1 _1152_ (.A1(\current_multiplier[3] ),
    .A2(net157),
    .B1(net153),
    .B2(\current_multiplier[2] ),
    .C1(_0830_),
    .X(_0366_));
 sky130_fd_sc_hd__or2_1 _1153_ (.A(net44),
    .B(net208),
    .X(_0831_));
 sky130_fd_sc_hd__o221a_1 _1154_ (.A1(\current_multiplier[2] ),
    .A2(net156),
    .B1(net152),
    .B2(\current_multiplier[1] ),
    .C1(_0831_),
    .X(_0365_));
 sky130_fd_sc_hd__or2_1 _1155_ (.A(net33),
    .B(net205),
    .X(_0832_));
 sky130_fd_sc_hd__o221a_1 _1156_ (.A1(\current_multiplier[1] ),
    .A2(net156),
    .B1(net152),
    .B2(\current_multiplier[0] ),
    .C1(_0832_),
    .X(_0364_));
 sky130_fd_sc_hd__or4_4 _1157_ (.A(\extended_operand[15] ),
    .B(\extended_operand[14] ),
    .C(\extended_operand[13] ),
    .D(\extended_operand[12] ),
    .X(_0833_));
 sky130_fd_sc_hd__or4_4 _1158_ (.A(\extended_operand[3] ),
    .B(\extended_operand[2] ),
    .C(\extended_operand[1] ),
    .D(\extended_operand[0] ),
    .X(_0834_));
 sky130_fd_sc_hd__or4_1 _1159_ (.A(\extended_operand[7] ),
    .B(\extended_operand[6] ),
    .C(\extended_operand[5] ),
    .D(\extended_operand[4] ),
    .X(_0835_));
 sky130_fd_sc_hd__or4_1 _1160_ (.A(\extended_operand[11] ),
    .B(\extended_operand[10] ),
    .C(\extended_operand[9] ),
    .D(\extended_operand[8] ),
    .X(_0836_));
 sky130_fd_sc_hd__or3_2 _1161_ (.A(_0834_),
    .B(_0835_),
    .C(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__or3_1 _1162_ (.A(\extended_operand[18] ),
    .B(\extended_operand[17] ),
    .C(\extended_operand[16] ),
    .X(_0838_));
 sky130_fd_sc_hd__or4_1 _1163_ (.A(\extended_operand[19] ),
    .B(\extended_operand[18] ),
    .C(\extended_operand[17] ),
    .D(\extended_operand[16] ),
    .X(_0839_));
 sky130_fd_sc_hd__or2_1 _1164_ (.A(\extended_operand[21] ),
    .B(\extended_operand[20] ),
    .X(_0840_));
 sky130_fd_sc_hd__or4_1 _1165_ (.A(\extended_operand[23] ),
    .B(\extended_operand[22] ),
    .C(_0839_),
    .D(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__or2_1 _1166_ (.A(\extended_operand[25] ),
    .B(\extended_operand[24] ),
    .X(_0842_));
 sky130_fd_sc_hd__or4_4 _1167_ (.A(_0833_),
    .B(net149),
    .C(_0841_),
    .D(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__or2_1 _1168_ (.A(\extended_operand[27] ),
    .B(\extended_operand[26] ),
    .X(_0844_));
 sky130_fd_sc_hd__or3_1 _1169_ (.A(\extended_operand[30] ),
    .B(\extended_operand[29] ),
    .C(\extended_operand[28] ),
    .X(_0845_));
 sky130_fd_sc_hd__nor3_1 _1170_ (.A(_0843_),
    .B(_0844_),
    .C(_0845_),
    .Y(_0846_));
 sky130_fd_sc_hd__and2b_1 _1171_ (.A_N(net212),
    .B(\current_state[1] ),
    .X(_0847_));
 sky130_fd_sc_hd__nand2b_1 _1172_ (.A_N(net212),
    .B(\current_state[1] ),
    .Y(_0848_));
 sky130_fd_sc_hd__nand3b_1 _1173_ (.A_N(net212),
    .B(\current_state[0] ),
    .C(\current_state[1] ),
    .Y(_0849_));
 sky130_fd_sc_hd__nand2_1 _1174_ (.A(_0782_),
    .B(net185),
    .Y(_0850_));
 sky130_fd_sc_hd__or2_1 _1175_ (.A(_0782_),
    .B(net185),
    .X(_0851_));
 sky130_fd_sc_hd__o21a_1 _1176_ (.A1(_0846_),
    .A2(_0850_),
    .B1(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__nand2_1 _1177_ (.A(\partial_sum[61] ),
    .B(net137),
    .Y(_0853_));
 sky130_fd_sc_hd__or2_1 _1178_ (.A(\partial_sum[61] ),
    .B(net137),
    .X(_0854_));
 sky130_fd_sc_hd__nand2_1 _1179_ (.A(_0853_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__nand2_1 _1180_ (.A(\partial_sum[60] ),
    .B(net138),
    .Y(_0856_));
 sky130_fd_sc_hd__or2_1 _1181_ (.A(\partial_sum[60] ),
    .B(net138),
    .X(_0857_));
 sky130_fd_sc_hd__nand2_1 _1182_ (.A(_0856_),
    .B(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__and2_1 _1183_ (.A(\partial_sum[53] ),
    .B(net136),
    .X(_0859_));
 sky130_fd_sc_hd__nor2_1 _1184_ (.A(\partial_sum[53] ),
    .B(net140),
    .Y(_0860_));
 sky130_fd_sc_hd__or2_1 _1185_ (.A(_0859_),
    .B(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__nand2_1 _1186_ (.A(\partial_sum[54] ),
    .B(net138),
    .Y(_0862_));
 sky130_fd_sc_hd__or2_1 _1187_ (.A(\partial_sum[54] ),
    .B(net138),
    .X(_0863_));
 sky130_fd_sc_hd__nand2_1 _1188_ (.A(_0862_),
    .B(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__nand2_1 _1189_ (.A(\partial_sum[55] ),
    .B(net138),
    .Y(_0865_));
 sky130_fd_sc_hd__or2_1 _1190_ (.A(\partial_sum[55] ),
    .B(net138),
    .X(_0866_));
 sky130_fd_sc_hd__nand2_1 _1191_ (.A(_0865_),
    .B(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__xor2_1 _1192_ (.A(\partial_sum[52] ),
    .B(net137),
    .X(_0868_));
 sky130_fd_sc_hd__or4b_1 _1193_ (.A(_0861_),
    .B(_0864_),
    .C(_0867_),
    .D_N(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__nand2_1 _1194_ (.A(\partial_sum[49] ),
    .B(_0852_),
    .Y(_0870_));
 sky130_fd_sc_hd__or2_1 _1195_ (.A(\partial_sum[49] ),
    .B(_0852_),
    .X(_0871_));
 sky130_fd_sc_hd__nand2_1 _1196_ (.A(_0870_),
    .B(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__nand2_1 _1197_ (.A(\partial_sum[48] ),
    .B(net137),
    .Y(_0873_));
 sky130_fd_sc_hd__or2_1 _1198_ (.A(\partial_sum[48] ),
    .B(net136),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_1 _1199_ (.A(_0873_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__nand2_1 _1200_ (.A(\partial_sum[50] ),
    .B(net137),
    .Y(_0876_));
 sky130_fd_sc_hd__or2_1 _1201_ (.A(\partial_sum[50] ),
    .B(net137),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_1 _1202_ (.A(_0876_),
    .B(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__xnor2_1 _1203_ (.A(\partial_sum[51] ),
    .B(net137),
    .Y(_0879_));
 sky130_fd_sc_hd__or4_1 _1204_ (.A(_0872_),
    .B(_0875_),
    .C(_0878_),
    .D(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__o31a_1 _1205_ (.A1(_0833_),
    .A2(net149),
    .A3(_0838_),
    .B1(net184),
    .X(_0881_));
 sky130_fd_sc_hd__xnor2_1 _1206_ (.A(\extended_operand[19] ),
    .B(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__nor2_1 _1207_ (.A(\partial_sum[19] ),
    .B(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__nand2_1 _1208_ (.A(\partial_sum[19] ),
    .B(_0882_),
    .Y(_0884_));
 sky130_fd_sc_hd__nand2b_1 _1209_ (.A_N(_0883_),
    .B(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__o21a_1 _1210_ (.A1(_0833_),
    .A2(net149),
    .B1(net184),
    .X(_0886_));
 sky130_fd_sc_hd__o31a_1 _1211_ (.A1(\extended_operand[16] ),
    .A2(_0833_),
    .A3(net149),
    .B1(net184),
    .X(_0887_));
 sky130_fd_sc_hd__or4_1 _1212_ (.A(\extended_operand[17] ),
    .B(\extended_operand[16] ),
    .C(_0833_),
    .D(net149),
    .X(_0888_));
 sky130_fd_sc_hd__a21oi_1 _1213_ (.A1(net184),
    .A2(_0888_),
    .B1(_0783_),
    .Y(_0889_));
 sky130_fd_sc_hd__and3_1 _1214_ (.A(_0783_),
    .B(net184),
    .C(_0888_),
    .X(_0890_));
 sky130_fd_sc_hd__or2_1 _1215_ (.A(_0889_),
    .B(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__or3_1 _1216_ (.A(_0777_),
    .B(_0889_),
    .C(_0890_),
    .X(_0892_));
 sky130_fd_sc_hd__xnor2_1 _1217_ (.A(_0777_),
    .B(_0891_),
    .Y(_0893_));
 sky130_fd_sc_hd__xnor2_1 _1218_ (.A(\extended_operand[16] ),
    .B(_0886_),
    .Y(_0894_));
 sky130_fd_sc_hd__nand2_1 _1219_ (.A(\partial_sum[16] ),
    .B(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__or2_1 _1220_ (.A(\partial_sum[16] ),
    .B(_0894_),
    .X(_0896_));
 sky130_fd_sc_hd__nand2_1 _1221_ (.A(_0895_),
    .B(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__xnor2_1 _1222_ (.A(\extended_operand[17] ),
    .B(_0887_),
    .Y(_0898_));
 sky130_fd_sc_hd__nor2_1 _1223_ (.A(\partial_sum[17] ),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_1 _1224_ (.A(\partial_sum[17] ),
    .B(_0898_),
    .Y(_0900_));
 sky130_fd_sc_hd__nand2b_1 _1225_ (.A_N(_0899_),
    .B(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__or4_1 _1226_ (.A(_0885_),
    .B(_0893_),
    .C(_0897_),
    .D(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__nand2_1 _1227_ (.A(net149),
    .B(net184),
    .Y(_0903_));
 sky130_fd_sc_hd__o31a_1 _1228_ (.A1(\extended_operand[13] ),
    .A2(\extended_operand[12] ),
    .A3(net149),
    .B1(net184),
    .X(_0904_));
 sky130_fd_sc_hd__o41a_1 _1229_ (.A1(\extended_operand[14] ),
    .A2(\extended_operand[13] ),
    .A3(\extended_operand[12] ),
    .A4(net149),
    .B1(net184),
    .X(_0905_));
 sky130_fd_sc_hd__xor2_1 _1230_ (.A(\extended_operand[15] ),
    .B(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__xnor2_1 _1231_ (.A(_0778_),
    .B(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__xor2_1 _1232_ (.A(\extended_operand[14] ),
    .B(_0904_),
    .X(_0908_));
 sky130_fd_sc_hd__nand2b_1 _1233_ (.A_N(_0908_),
    .B(\partial_sum[14] ),
    .Y(_0909_));
 sky130_fd_sc_hd__xnor2_1 _1234_ (.A(\partial_sum[14] ),
    .B(_0908_),
    .Y(_0910_));
 sky130_fd_sc_hd__nand2b_1 _1235_ (.A_N(_0907_),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__xor2_2 _1236_ (.A(\extended_operand[12] ),
    .B(_0903_),
    .X(_0912_));
 sky130_fd_sc_hd__xnor2_1 _1237_ (.A(\partial_sum[12] ),
    .B(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__o21a_1 _1238_ (.A1(\extended_operand[12] ),
    .A2(net149),
    .B1(net184),
    .X(_0914_));
 sky130_fd_sc_hd__xnor2_1 _1239_ (.A(\extended_operand[13] ),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__nor2_1 _1240_ (.A(\partial_sum[13] ),
    .B(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__and2_1 _1241_ (.A(\partial_sum[13] ),
    .B(_0915_),
    .X(_0917_));
 sky130_fd_sc_hd__nor2_1 _1242_ (.A(_0916_),
    .B(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__or3b_1 _1243_ (.A(_0911_),
    .B(_0913_),
    .C_N(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__o21a_1 _1244_ (.A1(_0834_),
    .A2(_0835_),
    .B1(net183),
    .X(_0920_));
 sky130_fd_sc_hd__o31a_1 _1245_ (.A1(\extended_operand[8] ),
    .A2(_0834_),
    .A3(_0835_),
    .B1(net183),
    .X(_0921_));
 sky130_fd_sc_hd__o21a_1 _1246_ (.A1(\extended_operand[10] ),
    .A2(\extended_operand[9] ),
    .B1(net183),
    .X(_0922_));
 sky130_fd_sc_hd__a21oi_1 _1247_ (.A1(\extended_operand[9] ),
    .A2(net183),
    .B1(_0921_),
    .Y(_0923_));
 sky130_fd_sc_hd__or2_1 _1248_ (.A(_0921_),
    .B(_0922_),
    .X(_0924_));
 sky130_fd_sc_hd__xnor2_1 _1249_ (.A(\extended_operand[11] ),
    .B(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__nor2_1 _1250_ (.A(\partial_sum[11] ),
    .B(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__nand2_1 _1251_ (.A(\partial_sum[11] ),
    .B(_0925_),
    .Y(_0927_));
 sky130_fd_sc_hd__xnor2_1 _1252_ (.A(\partial_sum[11] ),
    .B(_0925_),
    .Y(_0928_));
 sky130_fd_sc_hd__xnor2_1 _1253_ (.A(\extended_operand[10] ),
    .B(_0923_),
    .Y(_0929_));
 sky130_fd_sc_hd__xnor2_1 _1254_ (.A(_0779_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__xnor2_1 _1255_ (.A(\extended_operand[9] ),
    .B(_0921_),
    .Y(_0931_));
 sky130_fd_sc_hd__nor2_1 _1256_ (.A(\partial_sum[9] ),
    .B(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__nand2_1 _1257_ (.A(\partial_sum[9] ),
    .B(_0931_),
    .Y(_0933_));
 sky130_fd_sc_hd__xnor2_1 _1258_ (.A(\extended_operand[8] ),
    .B(_0920_),
    .Y(_0934_));
 sky130_fd_sc_hd__nand2_1 _1259_ (.A(\partial_sum[8] ),
    .B(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__o21a_1 _1260_ (.A1(_0932_),
    .A2(_0935_),
    .B1(_0933_),
    .X(_0936_));
 sky130_fd_sc_hd__o31a_1 _1261_ (.A1(_0928_),
    .A2(_0930_),
    .A3(_0936_),
    .B1(_0927_),
    .X(_0937_));
 sky130_fd_sc_hd__o31ai_1 _1262_ (.A1(_0779_),
    .A2(_0926_),
    .A3(_0929_),
    .B1(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__o31a_1 _1263_ (.A1(\extended_operand[2] ),
    .A2(\extended_operand[1] ),
    .A3(\extended_operand[0] ),
    .B1(net186),
    .X(_0939_));
 sky130_fd_sc_hd__xnor2_1 _1264_ (.A(\extended_operand[3] ),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__and2_1 _1265_ (.A(\partial_sum[3] ),
    .B(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__o21a_1 _1266_ (.A1(\extended_operand[1] ),
    .A2(\extended_operand[0] ),
    .B1(net186),
    .X(_0942_));
 sky130_fd_sc_hd__xnor2_1 _1267_ (.A(\extended_operand[2] ),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__and2_1 _1268_ (.A(\partial_sum[2] ),
    .B(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__and3_1 _1269_ (.A(\extended_operand[1] ),
    .B(\extended_operand[0] ),
    .C(net183),
    .X(_0945_));
 sky130_fd_sc_hd__a21oi_1 _1270_ (.A1(\extended_operand[0] ),
    .A2(net183),
    .B1(\extended_operand[1] ),
    .Y(_0946_));
 sky130_fd_sc_hd__o21a_1 _1271_ (.A1(_0945_),
    .A2(_0946_),
    .B1(\partial_sum[1] ),
    .X(_0947_));
 sky130_fd_sc_hd__or3_1 _1272_ (.A(\partial_sum[1] ),
    .B(_0945_),
    .C(_0946_),
    .X(_0948_));
 sky130_fd_sc_hd__and2b_1 _1273_ (.A_N(_0947_),
    .B(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__nand2b_1 _1274_ (.A_N(\partial_sum[0] ),
    .B(\extended_operand[0] ),
    .Y(_0950_));
 sky130_fd_sc_hd__a21o_1 _1275_ (.A1(_0948_),
    .A2(_0950_),
    .B1(_0947_),
    .X(_0951_));
 sky130_fd_sc_hd__or2_1 _1276_ (.A(\partial_sum[2] ),
    .B(_0943_),
    .X(_0952_));
 sky130_fd_sc_hd__nand2b_1 _1277_ (.A_N(_0944_),
    .B(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__a21o_1 _1278_ (.A1(_0951_),
    .A2(_0952_),
    .B1(_0944_),
    .X(_0954_));
 sky130_fd_sc_hd__nor2_1 _1279_ (.A(\partial_sum[3] ),
    .B(_0940_),
    .Y(_0955_));
 sky130_fd_sc_hd__nor2_1 _1280_ (.A(_0941_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__and2_1 _1281_ (.A(_0954_),
    .B(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__inv_2 _1282_ (.A(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__a21o_1 _1283_ (.A1(_0954_),
    .A2(_0956_),
    .B1(_0941_),
    .X(_0959_));
 sky130_fd_sc_hd__nand2_1 _1284_ (.A(_0834_),
    .B(net183),
    .Y(_0960_));
 sky130_fd_sc_hd__xor2_2 _1285_ (.A(\extended_operand[4] ),
    .B(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__xor2_1 _1286_ (.A(\partial_sum[4] ),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__nand2_1 _1287_ (.A(_0959_),
    .B(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__o21a_1 _1288_ (.A1(\extended_operand[4] ),
    .A2(_0834_),
    .B1(net183),
    .X(_0964_));
 sky130_fd_sc_hd__o41a_1 _1289_ (.A1(\extended_operand[6] ),
    .A2(\extended_operand[5] ),
    .A3(\extended_operand[4] ),
    .A4(_0834_),
    .B1(net183),
    .X(_0965_));
 sky130_fd_sc_hd__xnor2_1 _1290_ (.A(\extended_operand[7] ),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__or2_1 _1291_ (.A(\partial_sum[7] ),
    .B(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__xnor2_1 _1292_ (.A(\partial_sum[7] ),
    .B(_0966_),
    .Y(_0968_));
 sky130_fd_sc_hd__o31a_1 _1293_ (.A1(\extended_operand[5] ),
    .A2(\extended_operand[4] ),
    .A3(_0834_),
    .B1(net183),
    .X(_0969_));
 sky130_fd_sc_hd__xnor2_1 _1294_ (.A(\extended_operand[6] ),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__nand2_1 _1295_ (.A(\partial_sum[6] ),
    .B(_0970_),
    .Y(_0971_));
 sky130_fd_sc_hd__xnor2_1 _1296_ (.A(\partial_sum[6] ),
    .B(_0970_),
    .Y(_0972_));
 sky130_fd_sc_hd__nor2_1 _1297_ (.A(_0968_),
    .B(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__xnor2_1 _1298_ (.A(\extended_operand[5] ),
    .B(_0964_),
    .Y(_0974_));
 sky130_fd_sc_hd__nor2_1 _1299_ (.A(\partial_sum[5] ),
    .B(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__and2_1 _1300_ (.A(\partial_sum[5] ),
    .B(_0974_),
    .X(_0976_));
 sky130_fd_sc_hd__nor2_1 _1301_ (.A(_0975_),
    .B(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__and2_1 _1302_ (.A(_0962_),
    .B(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__a22oi_1 _1303_ (.A1(\partial_sum[4] ),
    .A2(_0961_),
    .B1(_0974_),
    .B2(\partial_sum[5] ),
    .Y(_0979_));
 sky130_fd_sc_hd__nor2_1 _1304_ (.A(_0975_),
    .B(_0979_),
    .Y(_0980_));
 sky130_fd_sc_hd__a22o_1 _1305_ (.A1(\partial_sum[7] ),
    .A2(_0966_),
    .B1(_0970_),
    .B2(\partial_sum[6] ),
    .X(_0981_));
 sky130_fd_sc_hd__a22o_1 _1306_ (.A1(_0973_),
    .A2(_0980_),
    .B1(_0981_),
    .B2(_0967_),
    .X(_0982_));
 sky130_fd_sc_hd__a31o_1 _1307_ (.A1(_0959_),
    .A2(_0973_),
    .A3(_0978_),
    .B1(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__nand2b_1 _1308_ (.A_N(_0932_),
    .B(_0933_),
    .Y(_0984_));
 sky130_fd_sc_hd__or2_1 _1309_ (.A(\partial_sum[8] ),
    .B(_0934_),
    .X(_0985_));
 sky130_fd_sc_hd__and2_1 _1310_ (.A(_0935_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__nor4b_1 _1311_ (.A(_0928_),
    .B(_0930_),
    .C(_0984_),
    .D_N(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__a21oi_1 _1312_ (.A1(_0983_),
    .A2(net132),
    .B1(_0938_),
    .Y(_0988_));
 sky130_fd_sc_hd__nand2b_1 _1313_ (.A_N(_0919_),
    .B(_0938_),
    .Y(_0989_));
 sky130_fd_sc_hd__nand3b_1 _1314_ (.A_N(_0919_),
    .B(_0983_),
    .C(net132),
    .Y(_0990_));
 sky130_fd_sc_hd__a22o_1 _1315_ (.A1(\partial_sum[12] ),
    .A2(_0912_),
    .B1(_0915_),
    .B2(\partial_sum[13] ),
    .X(_0991_));
 sky130_fd_sc_hd__or3b_1 _1316_ (.A(_0911_),
    .B(_0916_),
    .C_N(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__a21o_1 _1317_ (.A1(_0778_),
    .A2(_0906_),
    .B1(_0909_),
    .X(_0993_));
 sky130_fd_sc_hd__o211a_1 _1318_ (.A1(_0778_),
    .A2(_0906_),
    .B1(_0992_),
    .C1(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__and3_1 _1319_ (.A(_0989_),
    .B(_0990_),
    .C(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__a31o_2 _1320_ (.A1(_0989_),
    .A2(_0990_),
    .A3(_0994_),
    .B1(_0902_),
    .X(_0996_));
 sky130_fd_sc_hd__or4_1 _1321_ (.A(_0833_),
    .B(net149),
    .C(_0839_),
    .D(_0840_),
    .X(_0997_));
 sky130_fd_sc_hd__nand2_1 _1322_ (.A(net185),
    .B(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__o21ai_1 _1323_ (.A1(\extended_operand[22] ),
    .A2(_0997_),
    .B1(net185),
    .Y(_0999_));
 sky130_fd_sc_hd__xnor2_1 _1324_ (.A(\extended_operand[23] ),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__xnor2_1 _1325_ (.A(_0775_),
    .B(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__xnor2_1 _1326_ (.A(\extended_operand[22] ),
    .B(_0998_),
    .Y(_1002_));
 sky130_fd_sc_hd__xnor2_1 _1327_ (.A(_0776_),
    .B(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__o31a_1 _1328_ (.A1(_0833_),
    .A2(_0837_),
    .A3(_0839_),
    .B1(net184),
    .X(_1004_));
 sky130_fd_sc_hd__or4_1 _1329_ (.A(\extended_operand[20] ),
    .B(_0833_),
    .C(_0837_),
    .D(_0839_),
    .X(_1005_));
 sky130_fd_sc_hd__nand3b_1 _1330_ (.A_N(\extended_operand[21] ),
    .B(net185),
    .C(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__a21bo_1 _1331_ (.A1(net185),
    .A2(_1005_),
    .B1_N(\extended_operand[21] ),
    .X(_1007_));
 sky130_fd_sc_hd__a21oi_1 _1332_ (.A1(_1006_),
    .A2(_1007_),
    .B1(\partial_sum[21] ),
    .Y(_1008_));
 sky130_fd_sc_hd__xnor2_1 _1333_ (.A(\extended_operand[20] ),
    .B(_1004_),
    .Y(_1009_));
 sky130_fd_sc_hd__nand2_1 _1334_ (.A(\partial_sum[20] ),
    .B(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__or2_1 _1335_ (.A(\partial_sum[20] ),
    .B(_1009_),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_1 _1336_ (.A(_1010_),
    .B(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__nand3_1 _1337_ (.A(\partial_sum[21] ),
    .B(_1006_),
    .C(_1007_),
    .Y(_1013_));
 sky130_fd_sc_hd__nand2b_1 _1338_ (.A_N(_1008_),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__or4_2 _1339_ (.A(_1001_),
    .B(_1003_),
    .C(_1012_),
    .D(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__o31a_1 _1340_ (.A1(\extended_operand[28] ),
    .A2(_0843_),
    .A3(_0844_),
    .B1(net185),
    .X(_1016_));
 sky130_fd_sc_hd__o41a_1 _1341_ (.A1(\extended_operand[29] ),
    .A2(\extended_operand[28] ),
    .A3(_0843_),
    .A4(_0844_),
    .B1(net185),
    .X(_1017_));
 sky130_fd_sc_hd__xor2_1 _1342_ (.A(\extended_operand[30] ),
    .B(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__nand2b_1 _1343_ (.A_N(_1018_),
    .B(\partial_sum[30] ),
    .Y(_1019_));
 sky130_fd_sc_hd__xor2_1 _1344_ (.A(\partial_sum[30] ),
    .B(_1018_),
    .X(_1020_));
 sky130_fd_sc_hd__or4_1 _1345_ (.A(_0782_),
    .B(_0843_),
    .C(_0844_),
    .D(_0845_),
    .X(_1021_));
 sky130_fd_sc_hd__o211a_1 _1346_ (.A1(_0846_),
    .A2(_0850_),
    .B1(_0851_),
    .C1(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__nand2_1 _1347_ (.A(\partial_sum[31] ),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__nor2_1 _1348_ (.A(\partial_sum[31] ),
    .B(_1022_),
    .Y(_1024_));
 sky130_fd_sc_hd__xnor2_1 _1349_ (.A(\partial_sum[31] ),
    .B(_1022_),
    .Y(_1025_));
 sky130_fd_sc_hd__xnor2_1 _1350_ (.A(\extended_operand[29] ),
    .B(_1016_),
    .Y(_1026_));
 sky130_fd_sc_hd__nor2_1 _1351_ (.A(\partial_sum[29] ),
    .B(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__nand2_1 _1352_ (.A(\partial_sum[29] ),
    .B(_1026_),
    .Y(_1028_));
 sky130_fd_sc_hd__xnor2_1 _1353_ (.A(\partial_sum[29] ),
    .B(_1026_),
    .Y(_1029_));
 sky130_fd_sc_hd__o21a_1 _1354_ (.A1(_0843_),
    .A2(_0844_),
    .B1(net185),
    .X(_1030_));
 sky130_fd_sc_hd__xnor2_1 _1355_ (.A(\extended_operand[28] ),
    .B(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__nand2_1 _1356_ (.A(\partial_sum[28] ),
    .B(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__xnor2_1 _1357_ (.A(\partial_sum[28] ),
    .B(_1031_),
    .Y(_1033_));
 sky130_fd_sc_hd__or4_1 _1358_ (.A(_1020_),
    .B(_1025_),
    .C(_1029_),
    .D(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__inv_2 _1359_ (.A(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__o31a_1 _1360_ (.A1(_0833_),
    .A2(_0837_),
    .A3(_0841_),
    .B1(net185),
    .X(_1036_));
 sky130_fd_sc_hd__xnor2_1 _1361_ (.A(\extended_operand[24] ),
    .B(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__xnor2_1 _1362_ (.A(\partial_sum[24] ),
    .B(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__nand2_1 _1363_ (.A(_0843_),
    .B(net186),
    .Y(_1039_));
 sky130_fd_sc_hd__o21ai_1 _1364_ (.A1(\extended_operand[26] ),
    .A2(_0843_),
    .B1(net186),
    .Y(_1040_));
 sky130_fd_sc_hd__xnor2_1 _1365_ (.A(\extended_operand[27] ),
    .B(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__nand2_1 _1366_ (.A(_0773_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__xnor2_1 _1367_ (.A(\partial_sum[27] ),
    .B(_1041_),
    .Y(_1043_));
 sky130_fd_sc_hd__xor2_2 _1368_ (.A(\extended_operand[26] ),
    .B(_1039_),
    .X(_1044_));
 sky130_fd_sc_hd__xor2_1 _1369_ (.A(\partial_sum[26] ),
    .B(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__a21o_1 _1370_ (.A1(\extended_operand[24] ),
    .A2(net186),
    .B1(_1036_),
    .X(_1046_));
 sky130_fd_sc_hd__xor2_1 _1371_ (.A(\extended_operand[25] ),
    .B(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__nand2_1 _1372_ (.A(_0774_),
    .B(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__xnor2_1 _1373_ (.A(\partial_sum[25] ),
    .B(_1047_),
    .Y(_1049_));
 sky130_fd_sc_hd__and3_1 _1374_ (.A(_1043_),
    .B(_1045_),
    .C(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__or3b_1 _1375_ (.A(_1034_),
    .B(_1038_),
    .C_N(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__o21a_1 _1376_ (.A1(_0895_),
    .A2(_0899_),
    .B1(_0900_),
    .X(_1052_));
 sky130_fd_sc_hd__a21o_1 _1377_ (.A1(_0884_),
    .A2(_0892_),
    .B1(_0883_),
    .X(_1053_));
 sky130_fd_sc_hd__o31a_1 _1378_ (.A1(_0885_),
    .A2(_0893_),
    .A3(_1052_),
    .B1(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__a211o_1 _1379_ (.A1(_0775_),
    .A2(_1000_),
    .B1(_1002_),
    .C1(_0776_),
    .X(_1055_));
 sky130_fd_sc_hd__o21a_1 _1380_ (.A1(_0775_),
    .A2(_1000_),
    .B1(_1055_),
    .X(_0403_));
 sky130_fd_sc_hd__and2_1 _1381_ (.A(_1010_),
    .B(_1013_),
    .X(_0404_));
 sky130_fd_sc_hd__or4_1 _1382_ (.A(_1001_),
    .B(_1003_),
    .C(_1008_),
    .D(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__o211a_1 _1383_ (.A1(_1015_),
    .A2(_1054_),
    .B1(_0403_),
    .C1(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__a21o_1 _1384_ (.A1(_1028_),
    .A2(_1032_),
    .B1(_1027_),
    .X(_0407_));
 sky130_fd_sc_hd__or3_1 _1385_ (.A(_1020_),
    .B(_1025_),
    .C(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__o211a_1 _1386_ (.A1(_1019_),
    .A2(_1024_),
    .B1(_0408_),
    .C1(_1023_),
    .X(_0409_));
 sky130_fd_sc_hd__a2bb2o_1 _1387_ (.A1_N(_0774_),
    .A2_N(_1047_),
    .B1(_1037_),
    .B2(\partial_sum[24] ),
    .X(_0410_));
 sky130_fd_sc_hd__and3_1 _1388_ (.A(_1043_),
    .B(_1045_),
    .C(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__a2bb2o_1 _1389_ (.A1_N(_0773_),
    .A2_N(_1041_),
    .B1(_1044_),
    .B2(\partial_sum[26] ),
    .X(_0412_));
 sky130_fd_sc_hd__a22o_1 _1390_ (.A1(_1048_),
    .A2(_0411_),
    .B1(_0412_),
    .B2(_1042_),
    .X(_0413_));
 sky130_fd_sc_hd__o2bb2a_1 _1391_ (.A1_N(_1035_),
    .A2_N(_0413_),
    .B1(_1051_),
    .B2(_0406_),
    .X(_0414_));
 sky130_fd_sc_hd__o311ai_4 _1392_ (.A1(_0996_),
    .A2(_1015_),
    .A3(_1051_),
    .B1(_0409_),
    .C1(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__nand2_1 _1393_ (.A(\partial_sum[33] ),
    .B(net135),
    .Y(_0416_));
 sky130_fd_sc_hd__or2_1 _1394_ (.A(\partial_sum[33] ),
    .B(net135),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _1395_ (.A(_0416_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__xnor2_1 _1396_ (.A(\partial_sum[35] ),
    .B(net135),
    .Y(_0419_));
 sky130_fd_sc_hd__nand2_1 _1397_ (.A(\partial_sum[34] ),
    .B(net135),
    .Y(_0420_));
 sky130_fd_sc_hd__or2_1 _1398_ (.A(\partial_sum[34] ),
    .B(net135),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_1 _1399_ (.A(_0420_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__xnor2_1 _1400_ (.A(\partial_sum[32] ),
    .B(net135),
    .Y(_0423_));
 sky130_fd_sc_hd__or4_1 _1401_ (.A(_0418_),
    .B(_0419_),
    .C(_0422_),
    .D(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__nand2_1 _1402_ (.A(\partial_sum[36] ),
    .B(net136),
    .Y(_0425_));
 sky130_fd_sc_hd__or2_1 _1403_ (.A(\partial_sum[36] ),
    .B(net136),
    .X(_0426_));
 sky130_fd_sc_hd__and2_1 _1404_ (.A(_0425_),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _1405_ (.A(_0425_),
    .B(_0426_),
    .Y(_0428_));
 sky130_fd_sc_hd__and2_1 _1406_ (.A(\partial_sum[37] ),
    .B(net136),
    .X(_0429_));
 sky130_fd_sc_hd__nor2_1 _1407_ (.A(\partial_sum[37] ),
    .B(net136),
    .Y(_0430_));
 sky130_fd_sc_hd__or2_1 _1408_ (.A(_0429_),
    .B(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__xnor2_1 _1409_ (.A(\partial_sum[39] ),
    .B(net134),
    .Y(_0432_));
 sky130_fd_sc_hd__nand2_1 _1410_ (.A(\partial_sum[38] ),
    .B(net136),
    .Y(_0433_));
 sky130_fd_sc_hd__or2_1 _1411_ (.A(\partial_sum[38] ),
    .B(net136),
    .X(_0434_));
 sky130_fd_sc_hd__nand2_1 _1412_ (.A(_0433_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__or4_1 _1413_ (.A(_0428_),
    .B(_0431_),
    .C(_0432_),
    .D(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__nor2_1 _1414_ (.A(_0424_),
    .B(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_1 _1415_ (.A(\partial_sum[41] ),
    .B(net133),
    .Y(_0438_));
 sky130_fd_sc_hd__or2_1 _1416_ (.A(\partial_sum[41] ),
    .B(net133),
    .X(_0439_));
 sky130_fd_sc_hd__nand2_1 _1417_ (.A(_0438_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__xnor2_1 _1418_ (.A(\partial_sum[43] ),
    .B(net133),
    .Y(_0441_));
 sky130_fd_sc_hd__nand2_1 _1419_ (.A(\partial_sum[42] ),
    .B(net133),
    .Y(_0442_));
 sky130_fd_sc_hd__or2_1 _1420_ (.A(\partial_sum[42] ),
    .B(net133),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _1421_ (.A(_0442_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _1422_ (.A(\partial_sum[40] ),
    .B(net133),
    .Y(_0445_));
 sky130_fd_sc_hd__or2_1 _1423_ (.A(\partial_sum[40] ),
    .B(net133),
    .X(_0446_));
 sky130_fd_sc_hd__nand2_1 _1424_ (.A(_0445_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__or4_1 _1425_ (.A(_0440_),
    .B(_0441_),
    .C(_0444_),
    .D(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__and2_1 _1426_ (.A(\partial_sum[44] ),
    .B(net134),
    .X(_0449_));
 sky130_fd_sc_hd__nor2_1 _1427_ (.A(\partial_sum[44] ),
    .B(net134),
    .Y(_0450_));
 sky130_fd_sc_hd__nor2_1 _1428_ (.A(_0449_),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__nand2_1 _1429_ (.A(\partial_sum[45] ),
    .B(net133),
    .Y(_0452_));
 sky130_fd_sc_hd__nor2_1 _1430_ (.A(\partial_sum[45] ),
    .B(net134),
    .Y(_0453_));
 sky130_fd_sc_hd__or2_1 _1431_ (.A(\partial_sum[45] ),
    .B(net133),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_1 _1432_ (.A(_0452_),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__xnor2_1 _1433_ (.A(\partial_sum[47] ),
    .B(net134),
    .Y(_0456_));
 sky130_fd_sc_hd__nand2_1 _1434_ (.A(\partial_sum[46] ),
    .B(net134),
    .Y(_0457_));
 sky130_fd_sc_hd__or2_1 _1435_ (.A(\partial_sum[46] ),
    .B(net134),
    .X(_0458_));
 sky130_fd_sc_hd__nand2_1 _1436_ (.A(_0457_),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__nor3_1 _1437_ (.A(_0455_),
    .B(_0456_),
    .C(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__and3b_1 _1438_ (.A_N(_0448_),
    .B(_0451_),
    .C(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__o41a_1 _1439_ (.A1(\partial_sum[35] ),
    .A2(\partial_sum[34] ),
    .A3(\partial_sum[33] ),
    .A4(\partial_sum[32] ),
    .B1(net135),
    .X(_0462_));
 sky130_fd_sc_hd__o41a_1 _1440_ (.A1(\partial_sum[39] ),
    .A2(\partial_sum[38] ),
    .A3(\partial_sum[37] ),
    .A4(\partial_sum[36] ),
    .B1(net136),
    .X(_0463_));
 sky130_fd_sc_hd__or2_1 _1441_ (.A(_0462_),
    .B(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__o41a_1 _1442_ (.A1(\partial_sum[43] ),
    .A2(\partial_sum[42] ),
    .A3(\partial_sum[41] ),
    .A4(\partial_sum[40] ),
    .B1(net133),
    .X(_0465_));
 sky130_fd_sc_hd__o41a_1 _1443_ (.A1(\partial_sum[47] ),
    .A2(\partial_sum[46] ),
    .A3(\partial_sum[45] ),
    .A4(\partial_sum[44] ),
    .B1(net134),
    .X(_0466_));
 sky130_fd_sc_hd__or3_1 _1444_ (.A(_0464_),
    .B(_0465_),
    .C(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__a31oi_2 _1445_ (.A1(_0415_),
    .A2(_0437_),
    .A3(_0461_),
    .B1(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__nor2_1 _1446_ (.A(_0880_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__o41a_1 _1447_ (.A1(\partial_sum[51] ),
    .A2(\partial_sum[50] ),
    .A3(\partial_sum[49] ),
    .A4(\partial_sum[48] ),
    .B1(net137),
    .X(_0470_));
 sky130_fd_sc_hd__inv_2 _1448_ (.A(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__o21ai_1 _1449_ (.A1(\partial_sum[53] ),
    .A2(\partial_sum[52] ),
    .B1(net135),
    .Y(_0472_));
 sky130_fd_sc_hd__and3_1 _1450_ (.A(_0862_),
    .B(_0865_),
    .C(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__o31a_1 _1451_ (.A1(_0869_),
    .A2(_0880_),
    .A3(_0468_),
    .B1(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__xnor2_1 _1452_ (.A(\partial_sum[59] ),
    .B(net138),
    .Y(_0475_));
 sky130_fd_sc_hd__xnor2_1 _1453_ (.A(\partial_sum[57] ),
    .B(net138),
    .Y(_0476_));
 sky130_fd_sc_hd__and2_1 _1454_ (.A(\partial_sum[58] ),
    .B(net139),
    .X(_0477_));
 sky130_fd_sc_hd__nor2_1 _1455_ (.A(\partial_sum[58] ),
    .B(net139),
    .Y(_0478_));
 sky130_fd_sc_hd__nor2_1 _1456_ (.A(_0477_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__xnor2_1 _1457_ (.A(\partial_sum[56] ),
    .B(net138),
    .Y(_0480_));
 sky130_fd_sc_hd__or4_1 _1458_ (.A(_0476_),
    .B(_0477_),
    .C(_0478_),
    .D(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__a211o_1 _1459_ (.A1(_0471_),
    .A2(_0474_),
    .B1(_0475_),
    .C1(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__o21a_1 _1460_ (.A1(\partial_sum[57] ),
    .A2(\partial_sum[56] ),
    .B1(net139),
    .X(_0483_));
 sky130_fd_sc_hd__a211oi_1 _1461_ (.A1(\partial_sum[59] ),
    .A2(net139),
    .B1(_0477_),
    .C1(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__a21o_1 _1462_ (.A1(_0482_),
    .A2(_0484_),
    .B1(_0858_),
    .X(_0485_));
 sky130_fd_sc_hd__a211o_1 _1463_ (.A1(_0482_),
    .A2(_0484_),
    .B1(_0855_),
    .C1(_0858_),
    .X(_0486_));
 sky130_fd_sc_hd__nand2_1 _1464_ (.A(\partial_sum[62] ),
    .B(net137),
    .Y(_0487_));
 sky130_fd_sc_hd__or2_1 _1465_ (.A(\partial_sum[62] ),
    .B(net137),
    .X(_0488_));
 sky130_fd_sc_hd__nand2_1 _1466_ (.A(_0487_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__nand4_1 _1467_ (.A(_0853_),
    .B(_0856_),
    .C(_0486_),
    .D(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__a31o_1 _1468_ (.A1(_0853_),
    .A2(_0856_),
    .A3(_0486_),
    .B1(_0489_),
    .X(_0491_));
 sky130_fd_sc_hd__and3_1 _1469_ (.A(net193),
    .B(_0490_),
    .C(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__nor2_1 _1470_ (.A(net151),
    .B(net191),
    .Y(_0493_));
 sky130_fd_sc_hd__nand2_1 _1471_ (.A(_0791_),
    .B(net189),
    .Y(_0494_));
 sky130_fd_sc_hd__and3_1 _1472_ (.A(\partial_sum[63] ),
    .B(net212),
    .C(_0784_),
    .X(_0495_));
 sky130_fd_sc_hd__a211o_1 _1473_ (.A1(\partial_sum[62] ),
    .A2(net148),
    .B1(_0495_),
    .C1(_0492_),
    .X(_0363_));
 sky130_fd_sc_hd__a21oi_1 _1474_ (.A1(_0856_),
    .A2(_0485_),
    .B1(_0855_),
    .Y(_0496_));
 sky130_fd_sc_hd__a31o_1 _1475_ (.A1(_0855_),
    .A2(_0856_),
    .A3(_0485_),
    .B1(net188),
    .X(_0497_));
 sky130_fd_sc_hd__nor2_1 _1476_ (.A(_0496_),
    .B(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__a221o_1 _1477_ (.A1(\partial_sum[62] ),
    .A2(net165),
    .B1(net147),
    .B2(\partial_sum[61] ),
    .C1(_0498_),
    .X(_0362_));
 sky130_fd_sc_hd__nand3_1 _1478_ (.A(_0858_),
    .B(_0482_),
    .C(_0484_),
    .Y(_0499_));
 sky130_fd_sc_hd__a22o_1 _1479_ (.A1(\partial_sum[61] ),
    .A2(net164),
    .B1(net147),
    .B2(\partial_sum[60] ),
    .X(_0500_));
 sky130_fd_sc_hd__a31o_1 _1480_ (.A1(net193),
    .A2(_0485_),
    .A3(_0499_),
    .B1(_0500_),
    .X(_0361_));
 sky130_fd_sc_hd__a21oi_2 _1481_ (.A1(_0471_),
    .A2(_0474_),
    .B1(_0480_),
    .Y(_0501_));
 sky130_fd_sc_hd__a21oi_1 _1482_ (.A1(\partial_sum[56] ),
    .A2(net138),
    .B1(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__o22a_1 _1483_ (.A1(\partial_sum[57] ),
    .A2(net139),
    .B1(_0483_),
    .B2(_0501_),
    .X(_0503_));
 sky130_fd_sc_hd__o221a_1 _1484_ (.A1(\partial_sum[57] ),
    .A2(net139),
    .B1(_0483_),
    .B2(_0501_),
    .C1(_0479_),
    .X(_0504_));
 sky130_fd_sc_hd__nor2_1 _1485_ (.A(_0477_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__xnor2_1 _1486_ (.A(_0475_),
    .B(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__a22oi_1 _1487_ (.A1(\partial_sum[60] ),
    .A2(net164),
    .B1(net147),
    .B2(\partial_sum[59] ),
    .Y(_0507_));
 sky130_fd_sc_hd__o21ai_1 _1488_ (.A1(net188),
    .A2(_0506_),
    .B1(_0507_),
    .Y(_0360_));
 sky130_fd_sc_hd__nor2_1 _1489_ (.A(net188),
    .B(_0504_),
    .Y(_0508_));
 sky130_fd_sc_hd__o21a_1 _1490_ (.A1(_0479_),
    .A2(_0503_),
    .B1(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__a221o_1 _1491_ (.A1(\partial_sum[59] ),
    .A2(net164),
    .B1(net147),
    .B2(\partial_sum[58] ),
    .C1(_0509_),
    .X(_0359_));
 sky130_fd_sc_hd__nand2_1 _1492_ (.A(_0476_),
    .B(_0502_),
    .Y(_0510_));
 sky130_fd_sc_hd__o21a_1 _1493_ (.A1(_0476_),
    .A2(_0502_),
    .B1(net193),
    .X(_0511_));
 sky130_fd_sc_hd__a22o_1 _1494_ (.A1(\partial_sum[58] ),
    .A2(net164),
    .B1(net148),
    .B2(\partial_sum[57] ),
    .X(_0512_));
 sky130_fd_sc_hd__a21o_1 _1495_ (.A1(_0510_),
    .A2(_0511_),
    .B1(_0512_),
    .X(_0358_));
 sky130_fd_sc_hd__and3_1 _1496_ (.A(_0471_),
    .B(_0474_),
    .C(_0480_),
    .X(_0513_));
 sky130_fd_sc_hd__a22oi_1 _1497_ (.A1(\partial_sum[57] ),
    .A2(net164),
    .B1(net147),
    .B2(\partial_sum[56] ),
    .Y(_0514_));
 sky130_fd_sc_hd__o31ai_1 _1498_ (.A1(net187),
    .A2(_0501_),
    .A3(_0513_),
    .B1(_0514_),
    .Y(_0357_));
 sky130_fd_sc_hd__o21ai_2 _1499_ (.A1(_0469_),
    .A2(_0470_),
    .B1(_0868_),
    .Y(_0515_));
 sky130_fd_sc_hd__a21bo_1 _1500_ (.A1(\partial_sum[52] ),
    .A2(net135),
    .B1_N(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__a21o_1 _1501_ (.A1(_0472_),
    .A2(_0515_),
    .B1(_0860_),
    .X(_0517_));
 sky130_fd_sc_hd__a211o_1 _1502_ (.A1(_0472_),
    .A2(_0515_),
    .B1(_0860_),
    .C1(_0864_),
    .X(_0518_));
 sky130_fd_sc_hd__a21oi_1 _1503_ (.A1(_0862_),
    .A2(_0518_),
    .B1(_0867_),
    .Y(_0519_));
 sky130_fd_sc_hd__a31o_1 _1504_ (.A1(_0862_),
    .A2(_0867_),
    .A3(_0518_),
    .B1(net188),
    .X(_0520_));
 sky130_fd_sc_hd__nor2_1 _1505_ (.A(_0519_),
    .B(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__a221o_1 _1506_ (.A1(\partial_sum[56] ),
    .A2(net164),
    .B1(net147),
    .B2(\partial_sum[55] ),
    .C1(_0521_),
    .X(_0356_));
 sky130_fd_sc_hd__nand2_1 _1507_ (.A(_0864_),
    .B(_0517_),
    .Y(_0522_));
 sky130_fd_sc_hd__a22o_1 _1508_ (.A1(\partial_sum[55] ),
    .A2(net164),
    .B1(net147),
    .B2(\partial_sum[54] ),
    .X(_0523_));
 sky130_fd_sc_hd__a31o_1 _1509_ (.A1(net193),
    .A2(_0518_),
    .A3(_0522_),
    .B1(_0523_),
    .X(_0355_));
 sky130_fd_sc_hd__xor2_1 _1510_ (.A(_0861_),
    .B(_0516_),
    .X(_0524_));
 sky130_fd_sc_hd__nor2_1 _1511_ (.A(net187),
    .B(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__a221o_1 _1512_ (.A1(\partial_sum[54] ),
    .A2(net164),
    .B1(net147),
    .B2(\partial_sum[53] ),
    .C1(_0525_),
    .X(_0354_));
 sky130_fd_sc_hd__or3_1 _1513_ (.A(_0868_),
    .B(_0469_),
    .C(_0470_),
    .X(_0526_));
 sky130_fd_sc_hd__a22o_1 _1514_ (.A1(\partial_sum[53] ),
    .A2(net164),
    .B1(net147),
    .B2(\partial_sum[52] ),
    .X(_0527_));
 sky130_fd_sc_hd__a31o_1 _1515_ (.A1(net193),
    .A2(_0515_),
    .A3(_0526_),
    .B1(_0527_),
    .X(_0353_));
 sky130_fd_sc_hd__or2_1 _1516_ (.A(_0875_),
    .B(_0468_),
    .X(_0528_));
 sky130_fd_sc_hd__a21bo_1 _1517_ (.A1(_0873_),
    .A2(_0528_),
    .B1_N(_0871_),
    .X(_0529_));
 sky130_fd_sc_hd__a21o_1 _1518_ (.A1(_0870_),
    .A2(_0529_),
    .B1(_0878_),
    .X(_0530_));
 sky130_fd_sc_hd__nand3_1 _1519_ (.A(_0876_),
    .B(_0879_),
    .C(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__a21o_1 _1520_ (.A1(_0876_),
    .A2(_0530_),
    .B1(_0879_),
    .X(_0532_));
 sky130_fd_sc_hd__a22o_1 _1521_ (.A1(\partial_sum[52] ),
    .A2(net164),
    .B1(net147),
    .B2(\partial_sum[51] ),
    .X(_0533_));
 sky130_fd_sc_hd__a31o_1 _1522_ (.A1(net193),
    .A2(_0531_),
    .A3(_0532_),
    .B1(_0533_),
    .X(_0352_));
 sky130_fd_sc_hd__nand3_1 _1523_ (.A(_0870_),
    .B(_0878_),
    .C(_0529_),
    .Y(_0534_));
 sky130_fd_sc_hd__a22o_1 _1524_ (.A1(\partial_sum[51] ),
    .A2(net165),
    .B1(net148),
    .B2(\partial_sum[50] ),
    .X(_0535_));
 sky130_fd_sc_hd__a31o_1 _1525_ (.A1(net193),
    .A2(_0530_),
    .A3(_0534_),
    .B1(_0535_),
    .X(_0351_));
 sky130_fd_sc_hd__a21o_1 _1526_ (.A1(_0873_),
    .A2(_0528_),
    .B1(_0872_),
    .X(_0536_));
 sky130_fd_sc_hd__nand3_1 _1527_ (.A(_0872_),
    .B(_0873_),
    .C(_0528_),
    .Y(_0537_));
 sky130_fd_sc_hd__a22o_1 _1528_ (.A1(\partial_sum[50] ),
    .A2(net165),
    .B1(net148),
    .B2(\partial_sum[49] ),
    .X(_0538_));
 sky130_fd_sc_hd__a31o_1 _1529_ (.A1(net193),
    .A2(_0536_),
    .A3(_0537_),
    .B1(_0538_),
    .X(_0350_));
 sky130_fd_sc_hd__nand2_1 _1530_ (.A(_0875_),
    .B(_0468_),
    .Y(_0539_));
 sky130_fd_sc_hd__a22o_1 _1531_ (.A1(\partial_sum[49] ),
    .A2(net165),
    .B1(net148),
    .B2(\partial_sum[48] ),
    .X(_0540_));
 sky130_fd_sc_hd__a31o_1 _1532_ (.A1(net193),
    .A2(_0528_),
    .A3(_0539_),
    .B1(_0540_),
    .X(_0349_));
 sky130_fd_sc_hd__a21oi_1 _1533_ (.A1(_0415_),
    .A2(_0437_),
    .B1(_0464_),
    .Y(_0541_));
 sky130_fd_sc_hd__o21bai_1 _1534_ (.A1(_0448_),
    .A2(_0541_),
    .B1_N(_0465_),
    .Y(_0542_));
 sky130_fd_sc_hd__a21oi_1 _1535_ (.A1(_0451_),
    .A2(_0542_),
    .B1(_0449_),
    .Y(_0543_));
 sky130_fd_sc_hd__a21o_1 _1536_ (.A1(_0452_),
    .A2(_0543_),
    .B1(_0453_),
    .X(_0544_));
 sky130_fd_sc_hd__o21ai_1 _1537_ (.A1(_0459_),
    .A2(_0544_),
    .B1(_0457_),
    .Y(_0545_));
 sky130_fd_sc_hd__xnor2_1 _1538_ (.A(_0456_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__a22o_1 _1539_ (.A1(\partial_sum[48] ),
    .A2(net165),
    .B1(net148),
    .B2(\partial_sum[47] ),
    .X(_0547_));
 sky130_fd_sc_hd__a21o_1 _1540_ (.A1(net192),
    .A2(_0546_),
    .B1(_0547_),
    .X(_0348_));
 sky130_fd_sc_hd__xnor2_1 _1541_ (.A(_0459_),
    .B(_0544_),
    .Y(_0548_));
 sky130_fd_sc_hd__nor2_1 _1542_ (.A(net188),
    .B(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__a221o_1 _1543_ (.A1(\partial_sum[47] ),
    .A2(net165),
    .B1(net148),
    .B2(\partial_sum[46] ),
    .C1(_0549_),
    .X(_0347_));
 sky130_fd_sc_hd__or2_1 _1544_ (.A(_0455_),
    .B(_0543_),
    .X(_0550_));
 sky130_fd_sc_hd__nand2_1 _1545_ (.A(_0455_),
    .B(_0543_),
    .Y(_0551_));
 sky130_fd_sc_hd__a22o_1 _1546_ (.A1(\partial_sum[46] ),
    .A2(net159),
    .B1(net143),
    .B2(\partial_sum[45] ),
    .X(_0552_));
 sky130_fd_sc_hd__a31o_1 _1547_ (.A1(net194),
    .A2(_0550_),
    .A3(_0551_),
    .B1(_0552_),
    .X(_0346_));
 sky130_fd_sc_hd__a21oi_1 _1548_ (.A1(_0451_),
    .A2(_0542_),
    .B1(net189),
    .Y(_0553_));
 sky130_fd_sc_hd__o21a_1 _1549_ (.A1(_0451_),
    .A2(_0542_),
    .B1(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__a221o_1 _1550_ (.A1(\partial_sum[45] ),
    .A2(net159),
    .B1(net143),
    .B2(\partial_sum[44] ),
    .C1(_0554_),
    .X(_0345_));
 sky130_fd_sc_hd__or2_1 _1551_ (.A(_0447_),
    .B(_0541_),
    .X(_0555_));
 sky130_fd_sc_hd__a21bo_1 _1552_ (.A1(_0445_),
    .A2(_0555_),
    .B1_N(_0439_),
    .X(_0556_));
 sky130_fd_sc_hd__a21o_1 _1553_ (.A1(_0438_),
    .A2(_0556_),
    .B1(_0444_),
    .X(_0557_));
 sky130_fd_sc_hd__a21o_1 _1554_ (.A1(_0442_),
    .A2(_0557_),
    .B1(_0441_),
    .X(_0558_));
 sky130_fd_sc_hd__nand3_1 _1555_ (.A(_0441_),
    .B(_0442_),
    .C(_0557_),
    .Y(_0559_));
 sky130_fd_sc_hd__a22o_1 _1556_ (.A1(\partial_sum[44] ),
    .A2(net159),
    .B1(net143),
    .B2(\partial_sum[43] ),
    .X(_0560_));
 sky130_fd_sc_hd__a31o_1 _1557_ (.A1(net190),
    .A2(_0558_),
    .A3(_0559_),
    .B1(_0560_),
    .X(_0344_));
 sky130_fd_sc_hd__nand3_1 _1558_ (.A(_0438_),
    .B(_0444_),
    .C(_0556_),
    .Y(_0561_));
 sky130_fd_sc_hd__a22o_1 _1559_ (.A1(\partial_sum[43] ),
    .A2(net159),
    .B1(net143),
    .B2(\partial_sum[42] ),
    .X(_0562_));
 sky130_fd_sc_hd__a31o_1 _1560_ (.A1(net191),
    .A2(_0557_),
    .A3(_0561_),
    .B1(_0562_),
    .X(_0343_));
 sky130_fd_sc_hd__a21o_1 _1561_ (.A1(_0445_),
    .A2(_0555_),
    .B1(_0440_),
    .X(_0563_));
 sky130_fd_sc_hd__nand3_1 _1562_ (.A(_0440_),
    .B(_0445_),
    .C(_0555_),
    .Y(_0564_));
 sky130_fd_sc_hd__a22o_1 _1563_ (.A1(\partial_sum[42] ),
    .A2(net159),
    .B1(net143),
    .B2(\partial_sum[41] ),
    .X(_0565_));
 sky130_fd_sc_hd__a31o_1 _1564_ (.A1(net191),
    .A2(_0563_),
    .A3(_0564_),
    .B1(_0565_),
    .X(_0342_));
 sky130_fd_sc_hd__nand2_1 _1565_ (.A(_0447_),
    .B(_0541_),
    .Y(_0566_));
 sky130_fd_sc_hd__a22o_1 _1566_ (.A1(\partial_sum[41] ),
    .A2(net159),
    .B1(net143),
    .B2(\partial_sum[40] ),
    .X(_0567_));
 sky130_fd_sc_hd__a31o_1 _1567_ (.A1(net192),
    .A2(_0555_),
    .A3(_0566_),
    .B1(_0567_),
    .X(_0341_));
 sky130_fd_sc_hd__and2b_1 _1568_ (.A_N(_0424_),
    .B(_0415_),
    .X(_0568_));
 sky130_fd_sc_hd__o21ai_2 _1569_ (.A1(_0462_),
    .A2(_0568_),
    .B1(_0427_),
    .Y(_0569_));
 sky130_fd_sc_hd__a21oi_1 _1570_ (.A1(_0425_),
    .A2(_0569_),
    .B1(_0430_),
    .Y(_0570_));
 sky130_fd_sc_hd__nor2_1 _1571_ (.A(_0429_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__o21ai_1 _1572_ (.A1(_0435_),
    .A2(_0571_),
    .B1(_0433_),
    .Y(_0572_));
 sky130_fd_sc_hd__xnor2_1 _1573_ (.A(_0432_),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__a22o_1 _1574_ (.A1(\partial_sum[40] ),
    .A2(net163),
    .B1(net146),
    .B2(\partial_sum[39] ),
    .X(_0574_));
 sky130_fd_sc_hd__a21o_1 _1575_ (.A1(net192),
    .A2(_0573_),
    .B1(_0574_),
    .X(_0340_));
 sky130_fd_sc_hd__xnor2_1 _1576_ (.A(_0435_),
    .B(_0571_),
    .Y(_0575_));
 sky130_fd_sc_hd__nor2_1 _1577_ (.A(net187),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__a221o_1 _1578_ (.A1(\partial_sum[39] ),
    .A2(net163),
    .B1(net146),
    .B2(\partial_sum[38] ),
    .C1(_0576_),
    .X(_0339_));
 sky130_fd_sc_hd__a21oi_1 _1579_ (.A1(_0425_),
    .A2(_0569_),
    .B1(_0431_),
    .Y(_0577_));
 sky130_fd_sc_hd__a31o_1 _1580_ (.A1(_0425_),
    .A2(_0431_),
    .A3(_0569_),
    .B1(net187),
    .X(_0578_));
 sky130_fd_sc_hd__nor2_1 _1581_ (.A(_0577_),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__a221o_1 _1582_ (.A1(\partial_sum[38] ),
    .A2(net163),
    .B1(net146),
    .B2(\partial_sum[37] ),
    .C1(_0579_),
    .X(_0338_));
 sky130_fd_sc_hd__or3_1 _1583_ (.A(_0427_),
    .B(_0462_),
    .C(_0568_),
    .X(_0580_));
 sky130_fd_sc_hd__a22o_1 _1584_ (.A1(\partial_sum[37] ),
    .A2(net162),
    .B1(net145),
    .B2(\partial_sum[36] ),
    .X(_0581_));
 sky130_fd_sc_hd__a31o_1 _1585_ (.A1(net192),
    .A2(_0569_),
    .A3(_0580_),
    .B1(_0581_),
    .X(_0337_));
 sky130_fd_sc_hd__and2b_1 _1586_ (.A_N(_0423_),
    .B(_0415_),
    .X(_0582_));
 sky130_fd_sc_hd__a21o_1 _1587_ (.A1(\partial_sum[32] ),
    .A2(net135),
    .B1(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__nand2_1 _1588_ (.A(_0417_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__a21o_1 _1589_ (.A1(_0416_),
    .A2(_0584_),
    .B1(_0422_),
    .X(_0585_));
 sky130_fd_sc_hd__a21o_1 _1590_ (.A1(_0420_),
    .A2(_0585_),
    .B1(_0419_),
    .X(_0586_));
 sky130_fd_sc_hd__nand3_1 _1591_ (.A(_0419_),
    .B(_0420_),
    .C(_0585_),
    .Y(_0587_));
 sky130_fd_sc_hd__a22o_1 _1592_ (.A1(\partial_sum[36] ),
    .A2(net162),
    .B1(net145),
    .B2(\partial_sum[35] ),
    .X(_0588_));
 sky130_fd_sc_hd__a31o_1 _1593_ (.A1(net192),
    .A2(_0586_),
    .A3(_0587_),
    .B1(_0588_),
    .X(_0336_));
 sky130_fd_sc_hd__nand3_1 _1594_ (.A(_0416_),
    .B(_0422_),
    .C(_0584_),
    .Y(_0589_));
 sky130_fd_sc_hd__a22o_1 _1595_ (.A1(\partial_sum[35] ),
    .A2(net162),
    .B1(net145),
    .B2(\partial_sum[34] ),
    .X(_0590_));
 sky130_fd_sc_hd__a31o_1 _1596_ (.A1(net192),
    .A2(_0585_),
    .A3(_0589_),
    .B1(_0590_),
    .X(_0335_));
 sky130_fd_sc_hd__xnor2_1 _1597_ (.A(_0418_),
    .B(_0583_),
    .Y(_0591_));
 sky130_fd_sc_hd__a22o_1 _1598_ (.A1(\partial_sum[34] ),
    .A2(net162),
    .B1(net145),
    .B2(\partial_sum[33] ),
    .X(_0592_));
 sky130_fd_sc_hd__a21o_1 _1599_ (.A1(net192),
    .A2(_0591_),
    .B1(_0592_),
    .X(_0334_));
 sky130_fd_sc_hd__and2b_1 _1600_ (.A_N(_0415_),
    .B(_0423_),
    .X(_0593_));
 sky130_fd_sc_hd__a22oi_1 _1601_ (.A1(\partial_sum[33] ),
    .A2(net162),
    .B1(net145),
    .B2(\partial_sum[32] ),
    .Y(_0594_));
 sky130_fd_sc_hd__o31ai_1 _1602_ (.A1(net187),
    .A2(_0582_),
    .A3(_0593_),
    .B1(_0594_),
    .Y(_0333_));
 sky130_fd_sc_hd__or2_1 _1603_ (.A(_0996_),
    .B(_1015_),
    .X(_0595_));
 sky130_fd_sc_hd__a21oi_2 _1604_ (.A1(_0406_),
    .A2(_0595_),
    .B1(_1038_),
    .Y(_0596_));
 sky130_fd_sc_hd__a21oi_1 _1605_ (.A1(_1050_),
    .A2(_0596_),
    .B1(_0413_),
    .Y(_0597_));
 sky130_fd_sc_hd__or2_1 _1606_ (.A(_1033_),
    .B(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__nand2_1 _1607_ (.A(_1032_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__a311o_1 _1608_ (.A1(_1028_),
    .A2(_1032_),
    .A3(_0598_),
    .B1(_1027_),
    .C1(_1020_),
    .X(_0600_));
 sky130_fd_sc_hd__nand2_1 _1609_ (.A(_1019_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__xnor2_1 _1610_ (.A(_1025_),
    .B(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__a22o_1 _1611_ (.A1(\partial_sum[32] ),
    .A2(net162),
    .B1(net145),
    .B2(\partial_sum[31] ),
    .X(_0603_));
 sky130_fd_sc_hd__a21o_1 _1612_ (.A1(net192),
    .A2(_0602_),
    .B1(_0603_),
    .X(_0332_));
 sky130_fd_sc_hd__o211ai_1 _1613_ (.A1(_1027_),
    .A2(_0598_),
    .B1(_0407_),
    .C1(_1020_),
    .Y(_0604_));
 sky130_fd_sc_hd__a22o_1 _1614_ (.A1(\partial_sum[31] ),
    .A2(net162),
    .B1(net145),
    .B2(\partial_sum[30] ),
    .X(_0605_));
 sky130_fd_sc_hd__a31o_1 _1615_ (.A1(net192),
    .A2(_0600_),
    .A3(_0604_),
    .B1(_0605_),
    .X(_0331_));
 sky130_fd_sc_hd__xor2_1 _1616_ (.A(_1029_),
    .B(_0599_),
    .X(_0606_));
 sky130_fd_sc_hd__nor2_1 _1617_ (.A(net187),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__a221o_1 _1618_ (.A1(\partial_sum[30] ),
    .A2(net162),
    .B1(net145),
    .B2(\partial_sum[29] ),
    .C1(_0607_),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _1619_ (.A(_1033_),
    .B(_0597_),
    .Y(_0608_));
 sky130_fd_sc_hd__a22o_1 _1620_ (.A1(\partial_sum[29] ),
    .A2(net162),
    .B1(net145),
    .B2(\partial_sum[28] ),
    .X(_0609_));
 sky130_fd_sc_hd__a31o_1 _1621_ (.A1(net192),
    .A2(_0598_),
    .A3(_0608_),
    .B1(_0609_),
    .X(_0329_));
 sky130_fd_sc_hd__o21a_1 _1622_ (.A1(_0410_),
    .A2(_0596_),
    .B1(_1048_),
    .X(_0610_));
 sky130_fd_sc_hd__and2_1 _1623_ (.A(_1045_),
    .B(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__a21o_1 _1624_ (.A1(\partial_sum[26] ),
    .A2(_1044_),
    .B1(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__a21oi_1 _1625_ (.A1(_1043_),
    .A2(_0612_),
    .B1(net187),
    .Y(_0613_));
 sky130_fd_sc_hd__o21a_1 _1626_ (.A1(_1043_),
    .A2(_0612_),
    .B1(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__a221o_1 _1627_ (.A1(\partial_sum[28] ),
    .A2(net162),
    .B1(net145),
    .B2(\partial_sum[27] ),
    .C1(_0614_),
    .X(_0328_));
 sky130_fd_sc_hd__nor2_1 _1628_ (.A(_1045_),
    .B(_0610_),
    .Y(_0615_));
 sky130_fd_sc_hd__a22oi_1 _1629_ (.A1(\partial_sum[27] ),
    .A2(net163),
    .B1(net146),
    .B2(\partial_sum[26] ),
    .Y(_0616_));
 sky130_fd_sc_hd__o31ai_1 _1630_ (.A1(net187),
    .A2(_0611_),
    .A3(_0615_),
    .B1(_0616_),
    .Y(_0327_));
 sky130_fd_sc_hd__a21o_1 _1631_ (.A1(\partial_sum[24] ),
    .A2(_1037_),
    .B1(_0596_),
    .X(_0617_));
 sky130_fd_sc_hd__a21oi_1 _1632_ (.A1(_1049_),
    .A2(_0617_),
    .B1(net187),
    .Y(_0618_));
 sky130_fd_sc_hd__o21a_1 _1633_ (.A1(_1049_),
    .A2(_0617_),
    .B1(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__a221o_1 _1634_ (.A1(\partial_sum[26] ),
    .A2(net163),
    .B1(net146),
    .B2(\partial_sum[25] ),
    .C1(_0619_),
    .X(_0326_));
 sky130_fd_sc_hd__and3_1 _1635_ (.A(_1038_),
    .B(_0406_),
    .C(_0595_),
    .X(_0620_));
 sky130_fd_sc_hd__a22oi_1 _1636_ (.A1(\partial_sum[25] ),
    .A2(net163),
    .B1(net146),
    .B2(\partial_sum[24] ),
    .Y(_0621_));
 sky130_fd_sc_hd__o31ai_1 _1637_ (.A1(net187),
    .A2(_0596_),
    .A3(_0620_),
    .B1(_0621_),
    .Y(_0325_));
 sky130_fd_sc_hd__a21o_1 _1638_ (.A1(_0996_),
    .A2(_1054_),
    .B1(_1012_),
    .X(_0622_));
 sky130_fd_sc_hd__a21o_1 _1639_ (.A1(_0404_),
    .A2(_0622_),
    .B1(_1008_),
    .X(_0623_));
 sky130_fd_sc_hd__or2_1 _1640_ (.A(_1003_),
    .B(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__o21a_1 _1641_ (.A1(_0776_),
    .A2(_1002_),
    .B1(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__o21ai_1 _1642_ (.A1(_1001_),
    .A2(_0625_),
    .B1(net190),
    .Y(_0626_));
 sky130_fd_sc_hd__a21oi_1 _1643_ (.A1(_1001_),
    .A2(_0625_),
    .B1(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__a221o_1 _1644_ (.A1(\partial_sum[24] ),
    .A2(net163),
    .B1(net146),
    .B2(\partial_sum[23] ),
    .C1(_0627_),
    .X(_0324_));
 sky130_fd_sc_hd__nand2_1 _1645_ (.A(_1003_),
    .B(_0623_),
    .Y(_0628_));
 sky130_fd_sc_hd__a22o_1 _1646_ (.A1(\partial_sum[23] ),
    .A2(net159),
    .B1(net143),
    .B2(\partial_sum[22] ),
    .X(_0629_));
 sky130_fd_sc_hd__a31o_1 _1647_ (.A1(net191),
    .A2(_0624_),
    .A3(_0628_),
    .B1(_0629_),
    .X(_0323_));
 sky130_fd_sc_hd__a21oi_1 _1648_ (.A1(_1010_),
    .A2(_0622_),
    .B1(_1014_),
    .Y(_0630_));
 sky130_fd_sc_hd__a31o_1 _1649_ (.A1(_1010_),
    .A2(_1014_),
    .A3(_0622_),
    .B1(net189),
    .X(_0631_));
 sky130_fd_sc_hd__a22oi_1 _1650_ (.A1(\partial_sum[22] ),
    .A2(net159),
    .B1(net143),
    .B2(\partial_sum[21] ),
    .Y(_0632_));
 sky130_fd_sc_hd__o21ai_1 _1651_ (.A1(_0630_),
    .A2(_0631_),
    .B1(_0632_),
    .Y(_0322_));
 sky130_fd_sc_hd__nand3_1 _1652_ (.A(_0996_),
    .B(_1012_),
    .C(_1054_),
    .Y(_0633_));
 sky130_fd_sc_hd__a22o_1 _1653_ (.A1(\partial_sum[21] ),
    .A2(net159),
    .B1(net143),
    .B2(\partial_sum[20] ),
    .X(_0634_));
 sky130_fd_sc_hd__a31o_1 _1654_ (.A1(net191),
    .A2(_0622_),
    .A3(_0633_),
    .B1(_0634_),
    .X(_0321_));
 sky130_fd_sc_hd__or2_1 _1655_ (.A(_0897_),
    .B(_0995_),
    .X(_0635_));
 sky130_fd_sc_hd__a311o_1 _1656_ (.A1(_0895_),
    .A2(_0900_),
    .A3(_0635_),
    .B1(_0899_),
    .C1(_0893_),
    .X(_0636_));
 sky130_fd_sc_hd__nand3_1 _1657_ (.A(_0885_),
    .B(_0892_),
    .C(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__a21o_1 _1658_ (.A1(_0892_),
    .A2(_0636_),
    .B1(_0885_),
    .X(_0638_));
 sky130_fd_sc_hd__a22o_1 _1659_ (.A1(\partial_sum[20] ),
    .A2(net158),
    .B1(net142),
    .B2(\partial_sum[19] ),
    .X(_0639_));
 sky130_fd_sc_hd__a31o_1 _1660_ (.A1(net190),
    .A2(_0637_),
    .A3(_0638_),
    .B1(_0639_),
    .X(_0320_));
 sky130_fd_sc_hd__o211ai_1 _1661_ (.A1(_0901_),
    .A2(_0635_),
    .B1(_1052_),
    .C1(_0893_),
    .Y(_0640_));
 sky130_fd_sc_hd__a22o_1 _1662_ (.A1(\partial_sum[19] ),
    .A2(net158),
    .B1(net142),
    .B2(\partial_sum[18] ),
    .X(_0641_));
 sky130_fd_sc_hd__a31o_1 _1663_ (.A1(net190),
    .A2(_0636_),
    .A3(_0640_),
    .B1(_0641_),
    .X(_0319_));
 sky130_fd_sc_hd__nand3_1 _1664_ (.A(_0895_),
    .B(_0901_),
    .C(_0635_),
    .Y(_0642_));
 sky130_fd_sc_hd__a21o_1 _1665_ (.A1(_0895_),
    .A2(_0635_),
    .B1(_0901_),
    .X(_0643_));
 sky130_fd_sc_hd__a22o_1 _1666_ (.A1(\partial_sum[18] ),
    .A2(net158),
    .B1(net142),
    .B2(\partial_sum[17] ),
    .X(_0644_));
 sky130_fd_sc_hd__a31o_1 _1667_ (.A1(net190),
    .A2(_0642_),
    .A3(_0643_),
    .B1(_0644_),
    .X(_0318_));
 sky130_fd_sc_hd__nand2_1 _1668_ (.A(_0897_),
    .B(_0995_),
    .Y(_0645_));
 sky130_fd_sc_hd__a22o_1 _1669_ (.A1(\partial_sum[17] ),
    .A2(net158),
    .B1(net142),
    .B2(\partial_sum[16] ),
    .X(_0646_));
 sky130_fd_sc_hd__a31o_1 _1670_ (.A1(net190),
    .A2(_0635_),
    .A3(_0645_),
    .B1(_0646_),
    .X(_0317_));
 sky130_fd_sc_hd__nor2_1 _1671_ (.A(_0913_),
    .B(_0988_),
    .Y(_0647_));
 sky130_fd_sc_hd__nor2_1 _1672_ (.A(_0991_),
    .B(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__or3b_1 _1673_ (.A(_0916_),
    .B(_0648_),
    .C_N(_0910_),
    .X(_0649_));
 sky130_fd_sc_hd__a21oi_1 _1674_ (.A1(_0909_),
    .A2(_0649_),
    .B1(_0907_),
    .Y(_0650_));
 sky130_fd_sc_hd__a31o_1 _1675_ (.A1(_0907_),
    .A2(_0909_),
    .A3(_0649_),
    .B1(net189),
    .X(_0651_));
 sky130_fd_sc_hd__nor2_1 _1676_ (.A(_0650_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__a221o_1 _1677_ (.A1(\partial_sum[16] ),
    .A2(net158),
    .B1(net142),
    .B2(\partial_sum[15] ),
    .C1(_0652_),
    .X(_0316_));
 sky130_fd_sc_hd__o21ba_1 _1678_ (.A1(_0916_),
    .A2(_0648_),
    .B1_N(_0910_),
    .X(_0653_));
 sky130_fd_sc_hd__and3b_1 _1679_ (.A_N(_0653_),
    .B(net190),
    .C(_0649_),
    .X(_0654_));
 sky130_fd_sc_hd__a221o_1 _1680_ (.A1(\partial_sum[15] ),
    .A2(net158),
    .B1(net142),
    .B2(\partial_sum[14] ),
    .C1(_0654_),
    .X(_0315_));
 sky130_fd_sc_hd__a21o_1 _1681_ (.A1(\partial_sum[12] ),
    .A2(_0912_),
    .B1(_0647_),
    .X(_0655_));
 sky130_fd_sc_hd__a21oi_1 _1682_ (.A1(_0918_),
    .A2(_0655_),
    .B1(net189),
    .Y(_0656_));
 sky130_fd_sc_hd__o21a_1 _1683_ (.A1(_0918_),
    .A2(_0655_),
    .B1(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__a221o_1 _1684_ (.A1(\partial_sum[14] ),
    .A2(net158),
    .B1(net142),
    .B2(\partial_sum[13] ),
    .C1(_0657_),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _1685_ (.A(_0913_),
    .B(_0988_),
    .Y(_0658_));
 sky130_fd_sc_hd__and2b_1 _1686_ (.A_N(_0647_),
    .B(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__a221o_1 _1687_ (.A1(\partial_sum[13] ),
    .A2(net158),
    .B1(net190),
    .B2(_0659_),
    .C1(net142),
    .X(_0660_));
 sky130_fd_sc_hd__o21a_1 _1688_ (.A1(\partial_sum[12] ),
    .A2(net141),
    .B1(_0660_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _1689_ (.A(_0983_),
    .B(_0986_),
    .Y(_0661_));
 sky130_fd_sc_hd__a31o_1 _1690_ (.A1(_0933_),
    .A2(_0935_),
    .A3(_0661_),
    .B1(_0932_),
    .X(_0662_));
 sky130_fd_sc_hd__or2_1 _1691_ (.A(_0930_),
    .B(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__o21a_1 _1692_ (.A1(_0779_),
    .A2(_0929_),
    .B1(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__o21ai_1 _1693_ (.A1(_0928_),
    .A2(_0664_),
    .B1(net190),
    .Y(_0665_));
 sky130_fd_sc_hd__a21oi_1 _1694_ (.A1(_0928_),
    .A2(_0664_),
    .B1(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__a221o_1 _1695_ (.A1(\partial_sum[12] ),
    .A2(net158),
    .B1(net142),
    .B2(\partial_sum[11] ),
    .C1(_0666_),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_1 _1696_ (.A(_0930_),
    .B(_0662_),
    .Y(_0667_));
 sky130_fd_sc_hd__and3_1 _1697_ (.A(net190),
    .B(_0663_),
    .C(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__a21o_1 _1698_ (.A1(\partial_sum[11] ),
    .A2(net158),
    .B1(net142),
    .X(_0669_));
 sky130_fd_sc_hd__o22a_1 _1699_ (.A1(\partial_sum[10] ),
    .A2(net141),
    .B1(_0668_),
    .B2(_0669_),
    .X(_0311_));
 sky130_fd_sc_hd__nand2_1 _1700_ (.A(_0935_),
    .B(_0661_),
    .Y(_0670_));
 sky130_fd_sc_hd__xnor2_1 _1701_ (.A(_0984_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__a221o_1 _1702_ (.A1(\partial_sum[10] ),
    .A2(net160),
    .B1(net194),
    .B2(_0671_),
    .C1(net144),
    .X(_0672_));
 sky130_fd_sc_hd__o21a_1 _1703_ (.A1(\partial_sum[9] ),
    .A2(net141),
    .B1(_0672_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _1704_ (.A(_0983_),
    .B(_0986_),
    .X(_0673_));
 sky130_fd_sc_hd__a21o_1 _1705_ (.A1(\partial_sum[9] ),
    .A2(net160),
    .B1(net144),
    .X(_0674_));
 sky130_fd_sc_hd__a31o_1 _1706_ (.A1(net191),
    .A2(_0661_),
    .A3(_0673_),
    .B1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__o21a_1 _1707_ (.A1(\partial_sum[8] ),
    .A2(_0494_),
    .B1(_0675_),
    .X(_0309_));
 sky130_fd_sc_hd__a21bo_1 _1708_ (.A1(\partial_sum[4] ),
    .A2(_0961_),
    .B1_N(_0963_),
    .X(_0676_));
 sky130_fd_sc_hd__a21o_1 _1709_ (.A1(_0963_),
    .A2(_0979_),
    .B1(_0975_),
    .X(_0677_));
 sky130_fd_sc_hd__or2_1 _1710_ (.A(_0972_),
    .B(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__a21oi_1 _1711_ (.A1(_0971_),
    .A2(_0678_),
    .B1(_0968_),
    .Y(_0679_));
 sky130_fd_sc_hd__a31o_1 _1712_ (.A1(_0968_),
    .A2(_0971_),
    .A3(_0678_),
    .B1(net189),
    .X(_0680_));
 sky130_fd_sc_hd__nor2_1 _1713_ (.A(_0679_),
    .B(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__a21o_1 _1714_ (.A1(\partial_sum[8] ),
    .A2(net160),
    .B1(net144),
    .X(_0682_));
 sky130_fd_sc_hd__o22a_1 _1715_ (.A1(\partial_sum[7] ),
    .A2(net141),
    .B1(_0681_),
    .B2(_0682_),
    .X(_0308_));
 sky130_fd_sc_hd__nand2_1 _1716_ (.A(_0972_),
    .B(_0677_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _1717_ (.A(_0678_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__o221a_1 _1718_ (.A1(_0780_),
    .A2(net155),
    .B1(net189),
    .B2(_0684_),
    .C1(net141),
    .X(_0685_));
 sky130_fd_sc_hd__a21oi_1 _1719_ (.A1(_0781_),
    .A2(net144),
    .B1(_0685_),
    .Y(_0307_));
 sky130_fd_sc_hd__xnor2_1 _1720_ (.A(_0977_),
    .B(_0676_),
    .Y(_0686_));
 sky130_fd_sc_hd__o221a_1 _1721_ (.A1(_0781_),
    .A2(net155),
    .B1(net189),
    .B2(_0686_),
    .C1(net141),
    .X(_0687_));
 sky130_fd_sc_hd__o21ba_1 _1722_ (.A1(\partial_sum[5] ),
    .A2(net141),
    .B1_N(_0687_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _1723_ (.A(_0959_),
    .B(_0962_),
    .X(_0688_));
 sky130_fd_sc_hd__and3_1 _1724_ (.A(net194),
    .B(_0963_),
    .C(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__a21o_1 _1725_ (.A1(\partial_sum[5] ),
    .A2(net160),
    .B1(net144),
    .X(_0690_));
 sky130_fd_sc_hd__o22a_1 _1726_ (.A1(\partial_sum[4] ),
    .A2(_0494_),
    .B1(_0689_),
    .B2(_0690_),
    .X(_0305_));
 sky130_fd_sc_hd__or2_1 _1727_ (.A(_0954_),
    .B(_0956_),
    .X(_0691_));
 sky130_fd_sc_hd__a32o_1 _1728_ (.A1(net191),
    .A2(_0958_),
    .A3(_0691_),
    .B1(net160),
    .B2(\partial_sum[4] ),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _1729_ (.A0(\partial_sum[3] ),
    .A1(_0692_),
    .S(_0494_),
    .X(_0304_));
 sky130_fd_sc_hd__xnor2_1 _1730_ (.A(_0951_),
    .B(_0953_),
    .Y(_0693_));
 sky130_fd_sc_hd__a22o_1 _1731_ (.A1(\partial_sum[3] ),
    .A2(net160),
    .B1(net191),
    .B2(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _1732_ (.A0(\partial_sum[2] ),
    .A1(_0694_),
    .S(net141),
    .X(_0303_));
 sky130_fd_sc_hd__xor2_1 _1733_ (.A(_0949_),
    .B(_0950_),
    .X(_0695_));
 sky130_fd_sc_hd__a221o_1 _1734_ (.A1(\partial_sum[2] ),
    .A2(net161),
    .B1(net191),
    .B2(_0695_),
    .C1(net144),
    .X(_0696_));
 sky130_fd_sc_hd__o21a_1 _1735_ (.A1(\partial_sum[1] ),
    .A2(net141),
    .B1(_0696_),
    .X(_0302_));
 sky130_fd_sc_hd__o21ai_1 _1736_ (.A1(\extended_operand[0] ),
    .A2(net189),
    .B1(net141),
    .Y(_0697_));
 sky130_fd_sc_hd__a2bb2o_1 _1737_ (.A1_N(net189),
    .A2_N(_0950_),
    .B1(_0697_),
    .B2(\partial_sum[0] ),
    .X(_0698_));
 sky130_fd_sc_hd__a21o_1 _1738_ (.A1(\partial_sum[1] ),
    .A2(net161),
    .B1(_0698_),
    .X(_0301_));
 sky130_fd_sc_hd__and3b_1 _1739_ (.A_N(\current_state[1] ),
    .B(\current_state[0] ),
    .C(net212),
    .X(_0699_));
 sky130_fd_sc_hd__nand3b_2 _1740_ (.A_N(\current_state[1] ),
    .B(\current_state[0] ),
    .C(net212),
    .Y(_0700_));
 sky130_fd_sc_hd__a21o_1 _1741_ (.A1(net67),
    .A2(net203),
    .B1(net176),
    .X(_0300_));
 sky130_fd_sc_hd__and3_1 _1742_ (.A(net127),
    .B(net199),
    .C(net173),
    .X(_0701_));
 sky130_fd_sc_hd__a21o_1 _1743_ (.A1(\partial_sum[31] ),
    .A2(net181),
    .B1(_0701_),
    .X(_0299_));
 sky130_fd_sc_hd__and3_1 _1744_ (.A(net126),
    .B(net200),
    .C(net173),
    .X(_0702_));
 sky130_fd_sc_hd__a21o_1 _1745_ (.A1(\partial_sum[30] ),
    .A2(net181),
    .B1(_0702_),
    .X(_0298_));
 sky130_fd_sc_hd__and3_1 _1746_ (.A(net125),
    .B(net199),
    .C(net173),
    .X(_0703_));
 sky130_fd_sc_hd__a21o_1 _1747_ (.A1(\partial_sum[29] ),
    .A2(net181),
    .B1(_0703_),
    .X(_0297_));
 sky130_fd_sc_hd__and3_1 _1748_ (.A(net124),
    .B(net200),
    .C(net173),
    .X(_0704_));
 sky130_fd_sc_hd__a21o_1 _1749_ (.A1(\partial_sum[28] ),
    .A2(net181),
    .B1(_0704_),
    .X(_0296_));
 sky130_fd_sc_hd__and3_1 _1750_ (.A(net122),
    .B(net200),
    .C(net173),
    .X(_0705_));
 sky130_fd_sc_hd__a21o_1 _1751_ (.A1(\partial_sum[27] ),
    .A2(net181),
    .B1(_0705_),
    .X(_0295_));
 sky130_fd_sc_hd__and3_1 _1752_ (.A(net121),
    .B(net200),
    .C(net173),
    .X(_0706_));
 sky130_fd_sc_hd__a21o_1 _1753_ (.A1(\partial_sum[26] ),
    .A2(net181),
    .B1(_0706_),
    .X(_0294_));
 sky130_fd_sc_hd__and3_1 _1754_ (.A(net120),
    .B(net200),
    .C(net173),
    .X(_0707_));
 sky130_fd_sc_hd__a21o_1 _1755_ (.A1(\partial_sum[25] ),
    .A2(net181),
    .B1(_0707_),
    .X(_0293_));
 sky130_fd_sc_hd__and3_1 _1756_ (.A(net119),
    .B(net200),
    .C(net173),
    .X(_0708_));
 sky130_fd_sc_hd__a21o_1 _1757_ (.A1(\partial_sum[24] ),
    .A2(net181),
    .B1(_0708_),
    .X(_0292_));
 sky130_fd_sc_hd__and3_1 _1758_ (.A(net118),
    .B(net200),
    .C(net173),
    .X(_0709_));
 sky130_fd_sc_hd__a21o_1 _1759_ (.A1(\partial_sum[23] ),
    .A2(net181),
    .B1(_0709_),
    .X(_0291_));
 sky130_fd_sc_hd__and3_1 _1760_ (.A(net117),
    .B(net196),
    .C(net166),
    .X(_0710_));
 sky130_fd_sc_hd__a21o_1 _1761_ (.A1(\partial_sum[22] ),
    .A2(net179),
    .B1(_0710_),
    .X(_0290_));
 sky130_fd_sc_hd__and3_1 _1762_ (.A(net116),
    .B(net196),
    .C(net171),
    .X(_0711_));
 sky130_fd_sc_hd__a21o_1 _1763_ (.A1(\partial_sum[21] ),
    .A2(net179),
    .B1(_0711_),
    .X(_0289_));
 sky130_fd_sc_hd__and3_1 _1764_ (.A(net115),
    .B(net195),
    .C(net171),
    .X(_0712_));
 sky130_fd_sc_hd__a21o_1 _1765_ (.A1(\partial_sum[20] ),
    .A2(net175),
    .B1(_0712_),
    .X(_0288_));
 sky130_fd_sc_hd__and3_1 _1766_ (.A(net114),
    .B(net196),
    .C(net171),
    .X(_0713_));
 sky130_fd_sc_hd__a21o_1 _1767_ (.A1(\partial_sum[19] ),
    .A2(net179),
    .B1(_0713_),
    .X(_0287_));
 sky130_fd_sc_hd__and3_1 _1768_ (.A(net113),
    .B(net195),
    .C(net166),
    .X(_0714_));
 sky130_fd_sc_hd__a21o_1 _1769_ (.A1(\partial_sum[18] ),
    .A2(net175),
    .B1(_0714_),
    .X(_0286_));
 sky130_fd_sc_hd__and3_1 _1770_ (.A(net111),
    .B(net195),
    .C(net166),
    .X(_0715_));
 sky130_fd_sc_hd__a21o_1 _1771_ (.A1(\partial_sum[17] ),
    .A2(net175),
    .B1(_0715_),
    .X(_0285_));
 sky130_fd_sc_hd__and3_1 _1772_ (.A(net110),
    .B(net195),
    .C(net166),
    .X(_0716_));
 sky130_fd_sc_hd__a21o_1 _1773_ (.A1(\partial_sum[16] ),
    .A2(net175),
    .B1(_0716_),
    .X(_0284_));
 sky130_fd_sc_hd__and3_1 _1774_ (.A(net109),
    .B(net195),
    .C(net166),
    .X(_0717_));
 sky130_fd_sc_hd__a21o_1 _1775_ (.A1(\partial_sum[15] ),
    .A2(net175),
    .B1(_0717_),
    .X(_0283_));
 sky130_fd_sc_hd__and3_1 _1776_ (.A(net108),
    .B(net197),
    .C(net166),
    .X(_0718_));
 sky130_fd_sc_hd__a21o_1 _1777_ (.A1(\partial_sum[14] ),
    .A2(net175),
    .B1(_0718_),
    .X(_0282_));
 sky130_fd_sc_hd__and3_1 _1778_ (.A(net107),
    .B(net197),
    .C(net166),
    .X(_0719_));
 sky130_fd_sc_hd__a21o_1 _1779_ (.A1(\partial_sum[13] ),
    .A2(net175),
    .B1(_0719_),
    .X(_0281_));
 sky130_fd_sc_hd__and3_1 _1780_ (.A(net106),
    .B(net198),
    .C(net166),
    .X(_0720_));
 sky130_fd_sc_hd__a21o_1 _1781_ (.A1(\partial_sum[12] ),
    .A2(net175),
    .B1(_0720_),
    .X(_0280_));
 sky130_fd_sc_hd__and3_1 _1782_ (.A(net105),
    .B(net197),
    .C(net166),
    .X(_0721_));
 sky130_fd_sc_hd__a21o_1 _1783_ (.A1(\partial_sum[11] ),
    .A2(net175),
    .B1(_0721_),
    .X(_0279_));
 sky130_fd_sc_hd__and3_1 _1784_ (.A(net104),
    .B(net197),
    .C(net166),
    .X(_0722_));
 sky130_fd_sc_hd__a21o_1 _1785_ (.A1(\partial_sum[10] ),
    .A2(net175),
    .B1(_0722_),
    .X(_0278_));
 sky130_fd_sc_hd__and3_1 _1786_ (.A(net103),
    .B(net201),
    .C(net167),
    .X(_0723_));
 sky130_fd_sc_hd__a21o_1 _1787_ (.A1(\partial_sum[9] ),
    .A2(net177),
    .B1(_0723_),
    .X(_0277_));
 sky130_fd_sc_hd__and3_1 _1788_ (.A(net102),
    .B(net201),
    .C(net167),
    .X(_0724_));
 sky130_fd_sc_hd__a21o_1 _1789_ (.A1(\partial_sum[8] ),
    .A2(net177),
    .B1(_0724_),
    .X(_0276_));
 sky130_fd_sc_hd__and3_1 _1790_ (.A(net100),
    .B(net203),
    .C(net167),
    .X(_0725_));
 sky130_fd_sc_hd__a21o_1 _1791_ (.A1(\partial_sum[7] ),
    .A2(net176),
    .B1(_0725_),
    .X(_0275_));
 sky130_fd_sc_hd__and3_1 _1792_ (.A(net99),
    .B(net205),
    .C(net169),
    .X(_0726_));
 sky130_fd_sc_hd__a21o_1 _1793_ (.A1(\partial_sum[6] ),
    .A2(net178),
    .B1(_0726_),
    .X(_0274_));
 sky130_fd_sc_hd__and3_1 _1794_ (.A(net98),
    .B(net201),
    .C(net167),
    .X(_0727_));
 sky130_fd_sc_hd__a21o_1 _1795_ (.A1(\partial_sum[5] ),
    .A2(net177),
    .B1(_0727_),
    .X(_0273_));
 sky130_fd_sc_hd__and3_1 _1796_ (.A(net97),
    .B(net201),
    .C(net167),
    .X(_0728_));
 sky130_fd_sc_hd__a21o_1 _1797_ (.A1(\partial_sum[4] ),
    .A2(net177),
    .B1(_0728_),
    .X(_0272_));
 sky130_fd_sc_hd__and3_1 _1798_ (.A(net96),
    .B(net201),
    .C(net167),
    .X(_0729_));
 sky130_fd_sc_hd__a21o_1 _1799_ (.A1(\partial_sum[3] ),
    .A2(net177),
    .B1(_0729_),
    .X(_0271_));
 sky130_fd_sc_hd__and3_1 _1800_ (.A(net95),
    .B(net200),
    .C(net173),
    .X(_0730_));
 sky130_fd_sc_hd__a21o_1 _1801_ (.A1(\partial_sum[2] ),
    .A2(net181),
    .B1(_0730_),
    .X(_0270_));
 sky130_fd_sc_hd__and3_1 _1802_ (.A(net94),
    .B(net211),
    .C(net174),
    .X(_0731_));
 sky130_fd_sc_hd__a21o_1 _1803_ (.A1(\partial_sum[1] ),
    .A2(net182),
    .B1(_0731_),
    .X(_0269_));
 sky130_fd_sc_hd__and3_1 _1804_ (.A(net93),
    .B(net201),
    .C(net167),
    .X(_0732_));
 sky130_fd_sc_hd__a21o_1 _1805_ (.A1(\partial_sum[0] ),
    .A2(net177),
    .B1(_0732_),
    .X(_0268_));
 sky130_fd_sc_hd__and3_1 _1806_ (.A(net92),
    .B(net205),
    .C(net170),
    .X(_0733_));
 sky130_fd_sc_hd__a21o_1 _1807_ (.A1(\current_multiplier[31] ),
    .A2(net178),
    .B1(_0733_),
    .X(_0267_));
 sky130_fd_sc_hd__and3_1 _1808_ (.A(net91),
    .B(net205),
    .C(net170),
    .X(_0734_));
 sky130_fd_sc_hd__a21o_1 _1809_ (.A1(\current_multiplier[30] ),
    .A2(net178),
    .B1(_0734_),
    .X(_0266_));
 sky130_fd_sc_hd__and3_1 _1810_ (.A(net89),
    .B(net204),
    .C(net169),
    .X(_0735_));
 sky130_fd_sc_hd__a21o_1 _1811_ (.A1(\current_multiplier[29] ),
    .A2(net178),
    .B1(_0735_),
    .X(_0265_));
 sky130_fd_sc_hd__and3_1 _1812_ (.A(net88),
    .B(net205),
    .C(net169),
    .X(_0736_));
 sky130_fd_sc_hd__a21o_1 _1813_ (.A1(\current_multiplier[28] ),
    .A2(net178),
    .B1(_0736_),
    .X(_0264_));
 sky130_fd_sc_hd__and3_1 _1814_ (.A(net87),
    .B(net204),
    .C(net169),
    .X(_0737_));
 sky130_fd_sc_hd__a21o_1 _1815_ (.A1(\current_multiplier[27] ),
    .A2(net178),
    .B1(_0737_),
    .X(_0263_));
 sky130_fd_sc_hd__and3_1 _1816_ (.A(net86),
    .B(net204),
    .C(net169),
    .X(_0738_));
 sky130_fd_sc_hd__a21o_1 _1817_ (.A1(\current_multiplier[26] ),
    .A2(net178),
    .B1(_0738_),
    .X(_0262_));
 sky130_fd_sc_hd__and3_1 _1818_ (.A(net85),
    .B(net202),
    .C(net167),
    .X(_0739_));
 sky130_fd_sc_hd__a21o_1 _1819_ (.A1(\current_multiplier[25] ),
    .A2(net176),
    .B1(_0739_),
    .X(_0261_));
 sky130_fd_sc_hd__and3_1 _1820_ (.A(net84),
    .B(net203),
    .C(net167),
    .X(_0740_));
 sky130_fd_sc_hd__a21o_1 _1821_ (.A1(\current_multiplier[24] ),
    .A2(net176),
    .B1(_0740_),
    .X(_0260_));
 sky130_fd_sc_hd__and3_1 _1822_ (.A(net83),
    .B(net202),
    .C(net167),
    .X(_0741_));
 sky130_fd_sc_hd__a21o_1 _1823_ (.A1(\current_multiplier[23] ),
    .A2(net176),
    .B1(_0741_),
    .X(_0259_));
 sky130_fd_sc_hd__and3_1 _1824_ (.A(net82),
    .B(net202),
    .C(net168),
    .X(_0742_));
 sky130_fd_sc_hd__a21o_1 _1825_ (.A1(\current_multiplier[22] ),
    .A2(net176),
    .B1(_0742_),
    .X(_0258_));
 sky130_fd_sc_hd__and3_1 _1826_ (.A(net81),
    .B(net202),
    .C(net168),
    .X(_0743_));
 sky130_fd_sc_hd__a21o_1 _1827_ (.A1(\current_multiplier[21] ),
    .A2(net176),
    .B1(_0743_),
    .X(_0257_));
 sky130_fd_sc_hd__and3_1 _1828_ (.A(net80),
    .B(net203),
    .C(net168),
    .X(_0744_));
 sky130_fd_sc_hd__a21o_1 _1829_ (.A1(\current_multiplier[20] ),
    .A2(net176),
    .B1(_0744_),
    .X(_0256_));
 sky130_fd_sc_hd__and3_1 _1830_ (.A(net78),
    .B(net202),
    .C(net168),
    .X(_0745_));
 sky130_fd_sc_hd__a21o_1 _1831_ (.A1(\current_multiplier[19] ),
    .A2(net176),
    .B1(_0745_),
    .X(_0255_));
 sky130_fd_sc_hd__and3_1 _1832_ (.A(net77),
    .B(net205),
    .C(net169),
    .X(_0746_));
 sky130_fd_sc_hd__a21o_1 _1833_ (.A1(\current_multiplier[18] ),
    .A2(net177),
    .B1(_0746_),
    .X(_0254_));
 sky130_fd_sc_hd__and3_1 _1834_ (.A(net76),
    .B(net206),
    .C(net168),
    .X(_0747_));
 sky130_fd_sc_hd__a21o_1 _1835_ (.A1(\current_multiplier[17] ),
    .A2(net176),
    .B1(_0747_),
    .X(_0253_));
 sky130_fd_sc_hd__and3_1 _1836_ (.A(net75),
    .B(net204),
    .C(net169),
    .X(_0748_));
 sky130_fd_sc_hd__a21o_1 _1837_ (.A1(\current_multiplier[16] ),
    .A2(net178),
    .B1(_0748_),
    .X(_0252_));
 sky130_fd_sc_hd__and3_1 _1838_ (.A(net74),
    .B(net206),
    .C(net169),
    .X(_0749_));
 sky130_fd_sc_hd__a21o_1 _1839_ (.A1(\current_multiplier[15] ),
    .A2(net178),
    .B1(_0749_),
    .X(_0251_));
 sky130_fd_sc_hd__and3_1 _1840_ (.A(net73),
    .B(net204),
    .C(net169),
    .X(_0750_));
 sky130_fd_sc_hd__a21o_1 _1841_ (.A1(\current_multiplier[14] ),
    .A2(net179),
    .B1(_0750_),
    .X(_0250_));
 sky130_fd_sc_hd__and3_1 _1842_ (.A(net72),
    .B(net206),
    .C(net169),
    .X(_0751_));
 sky130_fd_sc_hd__a21o_1 _1843_ (.A1(\current_multiplier[13] ),
    .A2(net178),
    .B1(_0751_),
    .X(_0249_));
 sky130_fd_sc_hd__and3_1 _1844_ (.A(net71),
    .B(net208),
    .C(net172),
    .X(_0752_));
 sky130_fd_sc_hd__a21o_1 _1845_ (.A1(\current_multiplier[12] ),
    .A2(net180),
    .B1(_0752_),
    .X(_0248_));
 sky130_fd_sc_hd__and3_1 _1846_ (.A(net70),
    .B(net209),
    .C(net172),
    .X(_0753_));
 sky130_fd_sc_hd__a21o_1 _1847_ (.A1(\current_multiplier[11] ),
    .A2(net180),
    .B1(_0753_),
    .X(_0247_));
 sky130_fd_sc_hd__and3_1 _1848_ (.A(net69),
    .B(net209),
    .C(net172),
    .X(_0754_));
 sky130_fd_sc_hd__a21o_1 _1849_ (.A1(\current_multiplier[10] ),
    .A2(net180),
    .B1(_0754_),
    .X(_0246_));
 sky130_fd_sc_hd__and3_1 _1850_ (.A(net131),
    .B(net210),
    .C(net172),
    .X(_0755_));
 sky130_fd_sc_hd__a21o_1 _1851_ (.A1(\current_multiplier[9] ),
    .A2(net180),
    .B1(_0755_),
    .X(_0245_));
 sky130_fd_sc_hd__and3_1 _1852_ (.A(net130),
    .B(net210),
    .C(net172),
    .X(_0756_));
 sky130_fd_sc_hd__a21o_1 _1853_ (.A1(\current_multiplier[8] ),
    .A2(net180),
    .B1(_0756_),
    .X(_0244_));
 sky130_fd_sc_hd__and3_1 _1854_ (.A(net129),
    .B(net210),
    .C(net174),
    .X(_0757_));
 sky130_fd_sc_hd__a21o_1 _1855_ (.A1(\current_multiplier[7] ),
    .A2(net180),
    .B1(_0757_),
    .X(_0243_));
 sky130_fd_sc_hd__and3_1 _1856_ (.A(net128),
    .B(net210),
    .C(net172),
    .X(_0758_));
 sky130_fd_sc_hd__a21o_1 _1857_ (.A1(\current_multiplier[6] ),
    .A2(net182),
    .B1(_0758_),
    .X(_0242_));
 sky130_fd_sc_hd__and3_1 _1858_ (.A(net123),
    .B(net210),
    .C(net174),
    .X(_0759_));
 sky130_fd_sc_hd__a21o_1 _1859_ (.A1(\current_multiplier[5] ),
    .A2(net182),
    .B1(_0759_),
    .X(_0241_));
 sky130_fd_sc_hd__and3_1 _1860_ (.A(net112),
    .B(net210),
    .C(net174),
    .X(_0760_));
 sky130_fd_sc_hd__a21o_1 _1861_ (.A1(\current_multiplier[4] ),
    .A2(net182),
    .B1(_0760_),
    .X(_0240_));
 sky130_fd_sc_hd__and3_1 _1862_ (.A(net101),
    .B(net209),
    .C(net172),
    .X(_0761_));
 sky130_fd_sc_hd__a21o_1 _1863_ (.A1(\current_multiplier[3] ),
    .A2(net180),
    .B1(_0761_),
    .X(_0239_));
 sky130_fd_sc_hd__and3_1 _1864_ (.A(net90),
    .B(net208),
    .C(net172),
    .X(_0762_));
 sky130_fd_sc_hd__a21o_1 _1865_ (.A1(\current_multiplier[2] ),
    .A2(net180),
    .B1(_0762_),
    .X(_0238_));
 sky130_fd_sc_hd__and3_1 _1866_ (.A(net79),
    .B(net208),
    .C(net172),
    .X(_0763_));
 sky130_fd_sc_hd__a21o_1 _1867_ (.A1(\current_multiplier[1] ),
    .A2(net180),
    .B1(_0763_),
    .X(_0237_));
 sky130_fd_sc_hd__and3_1 _1868_ (.A(net68),
    .B(net209),
    .C(net172),
    .X(_0764_));
 sky130_fd_sc_hd__a21o_1 _1869_ (.A1(\current_multiplier[0] ),
    .A2(net180),
    .B1(_0764_),
    .X(_0236_));
 sky130_fd_sc_hd__xnor2_1 _1870_ (.A(\partial_sum[63] ),
    .B(net140),
    .Y(_0765_));
 sky130_fd_sc_hd__a21o_1 _1871_ (.A1(_0487_),
    .A2(_0491_),
    .B1(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__a31oi_1 _1872_ (.A1(_0487_),
    .A2(_0491_),
    .A3(_0765_),
    .B1(net188),
    .Y(_0767_));
 sky130_fd_sc_hd__a221o_1 _1873_ (.A1(\partial_sum[63] ),
    .A2(net148),
    .B1(_0766_),
    .B2(_0767_),
    .C1(_0495_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _1874_ (.A0(net25),
    .A1(\extended_operand[31] ),
    .S(net199),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _1875_ (.A0(net24),
    .A1(\extended_operand[30] ),
    .S(net199),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _1876_ (.A0(net22),
    .A1(\extended_operand[29] ),
    .S(net199),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _1877_ (.A0(net21),
    .A1(\extended_operand[28] ),
    .S(net199),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _1878_ (.A0(net20),
    .A1(\extended_operand[27] ),
    .S(net199),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _1879_ (.A0(net19),
    .A1(\extended_operand[26] ),
    .S(net199),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _1880_ (.A0(net18),
    .A1(\extended_operand[25] ),
    .S(net199),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _1881_ (.A0(net17),
    .A1(\extended_operand[24] ),
    .S(net199),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _1882_ (.A0(net16),
    .A1(\extended_operand[23] ),
    .S(net196),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _1883_ (.A0(net15),
    .A1(\extended_operand[22] ),
    .S(net196),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _1884_ (.A0(net14),
    .A1(\extended_operand[21] ),
    .S(net196),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _1885_ (.A0(net13),
    .A1(\extended_operand[20] ),
    .S(net196),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _1886_ (.A0(net11),
    .A1(\extended_operand[19] ),
    .S(net196),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _1887_ (.A0(net10),
    .A1(\extended_operand[18] ),
    .S(net195),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _1888_ (.A0(net9),
    .A1(\extended_operand[17] ),
    .S(net195),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _1889_ (.A0(net8),
    .A1(\extended_operand[16] ),
    .S(net195),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _1890_ (.A0(net7),
    .A1(\extended_operand[15] ),
    .S(net195),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _1891_ (.A0(net6),
    .A1(\extended_operand[14] ),
    .S(net195),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _1892_ (.A0(net5),
    .A1(\extended_operand[13] ),
    .S(net197),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _1893_ (.A0(net4),
    .A1(\extended_operand[12] ),
    .S(net197),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _1894_ (.A0(net3),
    .A1(\extended_operand[11] ),
    .S(net197),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _1895_ (.A0(net2),
    .A1(\extended_operand[10] ),
    .S(net197),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _1896_ (.A0(net32),
    .A1(\extended_operand[9] ),
    .S(net197),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _1897_ (.A0(net31),
    .A1(\extended_operand[8] ),
    .S(net201),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _1898_ (.A0(net30),
    .A1(\extended_operand[7] ),
    .S(net201),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _1899_ (.A0(net29),
    .A1(\extended_operand[6] ),
    .S(net207),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _1900_ (.A0(net28),
    .A1(\extended_operand[5] ),
    .S(net201),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _1901_ (.A0(net27),
    .A1(\extended_operand[4] ),
    .S(net201),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _1902_ (.A0(net26),
    .A1(\extended_operand[3] ),
    .S(net207),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _1903_ (.A0(net23),
    .A1(\extended_operand[2] ),
    .S(net197),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _1904_ (.A0(net12),
    .A1(\extended_operand[1] ),
    .S(net198),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _1905_ (.A0(net1),
    .A1(\extended_operand[0] ),
    .S(net198),
    .X(_0203_));
 sky130_fd_sc_hd__o21a_1 _1906_ (.A1(last_bit),
    .A2(_0772_),
    .B1(_0789_),
    .X(_0768_));
 sky130_fd_sc_hd__or3b_1 _1907_ (.A(net212),
    .B(\current_state[1] ),
    .C_N(\current_state[0] ),
    .X(_0769_));
 sky130_fd_sc_hd__o21ai_1 _1908_ (.A1(_0768_),
    .A2(_0769_),
    .B1(_0791_),
    .Y(\next_state[0] ));
 sky130_fd_sc_hd__xor2_1 _1909_ (.A(last_bit),
    .B(\current_multiplier[0] ),
    .X(_0770_));
 sky130_fd_sc_hd__and2_1 _1910_ (.A(_0789_),
    .B(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__and2b_1 _1911_ (.A_N(_0769_),
    .B(_0771_),
    .X(\next_state[1] ));
 sky130_fd_sc_hd__o21ai_1 _1912_ (.A1(_0769_),
    .A2(_0771_),
    .B1(net188),
    .Y(\next_state[2] ));
 sky130_fd_sc_hd__inv_2 _1913_ (.A(net217),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _1914_ (.A(net217),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1915_ (.A(net226),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _1916_ (.A(net225),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1917_ (.A(net225),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1918_ (.A(net225),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1919_ (.A(net225),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _1920_ (.A(net225),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1921_ (.A(net216),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1922_ (.A(net216),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _1923_ (.A(net216),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1924_ (.A(net216),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1925_ (.A(net216),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1926_ (.A(net213),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1927_ (.A(net213),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1928_ (.A(net213),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1929_ (.A(net213),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1930_ (.A(net213),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1931_ (.A(net213),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1932_ (.A(net214),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _1933_ (.A(net214),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1934_ (.A(net214),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1935_ (.A(net214),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1936_ (.A(net219),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1937_ (.A(net219),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1938_ (.A(net219),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1939_ (.A(net219),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1940_ (.A(net219),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1941_ (.A(net219),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1942_ (.A(net219),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _1943_ (.A(net219),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1944_ (.A(net234),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1945_ (.A(net230),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1946_ (.A(net231),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1947_ (.A(net236),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1948_ (.A(net236),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1949_ (.A(net236),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1950_ (.A(net238),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1951_ (.A(net238),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1952_ (.A(net238),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1953_ (.A(net238),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1954_ (.A(net238),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1955_ (.A(net237),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1956_ (.A(net237),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1957_ (.A(net237),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1958_ (.A(net231),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1959_ (.A(net231),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1960_ (.A(net231),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1961_ (.A(net231),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _1962_ (.A(net228),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _1963_ (.A(net229),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _1964_ (.A(net228),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _1965_ (.A(net229),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _1966_ (.A(net228),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _1967_ (.A(net228),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _1968_ (.A(net228),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _1969_ (.A(net228),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _1970_ (.A(net233),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _1971_ (.A(net231),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _1972_ (.A(net231),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _1973_ (.A(net230),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _1974_ (.A(net231),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _1975_ (.A(net230),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _1976_ (.A(net230),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _1977_ (.A(net225),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _1978_ (.A(net234),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _1979_ (.A(net221),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _1980_ (.A(net225),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _1981_ (.A(net227),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _1982_ (.A(net227),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _1983_ (.A(net230),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _1984_ (.A(net229),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _1985_ (.A(net225),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _1986_ (.A(net225),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1987_ (.A(net216),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _1988_ (.A(net216),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _1989_ (.A(net217),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _1990_ (.A(net216),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _1991_ (.A(net216),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _1992_ (.A(net213),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _1993_ (.A(net215),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _1994_ (.A(net213),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _1995_ (.A(net213),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _1996_ (.A(net214),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _1997_ (.A(net214),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _1998_ (.A(net214),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _1999_ (.A(net214),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _2000_ (.A(net221),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _2001_ (.A(net221),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _2002_ (.A(net221),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _2003_ (.A(net221),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _2004_ (.A(net223),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _2005_ (.A(net221),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _2006_ (.A(net219),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _2007_ (.A(net220),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _2008_ (.A(net220),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _2009_ (.A(net229),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _2010_ (.A(net226),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _2011_ (.A(net226),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _2012_ (.A(net226),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _2013_ (.A(net226),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _2014_ (.A(net226),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _2015_ (.A(net226),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _2016_ (.A(net230),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _2017_ (.A(net229),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _2018_ (.A(net225),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _2019_ (.A(net218),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _2020_ (.A(net218),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _2021_ (.A(net216),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _2022_ (.A(net217),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _2023_ (.A(net217),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _2024_ (.A(net217),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _2025_ (.A(net215),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _2026_ (.A(net215),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _2027_ (.A(net213),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _2028_ (.A(net214),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _2029_ (.A(net214),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _2030_ (.A(net215),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _2031_ (.A(net215),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _2032_ (.A(net217),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _2033_ (.A(net222),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _2034_ (.A(net219),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _2035_ (.A(net222),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _2036_ (.A(net222),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _2037_ (.A(net222),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _2038_ (.A(net220),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _2039_ (.A(net220),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _2040_ (.A(net220),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _2041_ (.A(net220),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _2042_ (.A(net221),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _2043_ (.A(net221),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _2044_ (.A(net221),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _2045_ (.A(net223),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _2046_ (.A(net221),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _2047_ (.A(net223),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _2048_ (.A(net222),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _2049_ (.A(net222),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _2050_ (.A(net222),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _2051_ (.A(net217),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _2052_ (.A(net217),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _2053_ (.A(net218),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _2054_ (.A(net218),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _2055_ (.A(net218),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _2056_ (.A(net234),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _2057_ (.A(net222),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _2058_ (.A(net222),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _2059_ (.A(net234),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _2060_ (.A(net234),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _2061_ (.A(net234),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _2062_ (.A(net222),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _2063_ (.A(net223),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _2064_ (.A(net235),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _2065_ (.A(net235),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _2066_ (.A(net235),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _2067_ (.A(net235),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _2068_ (.A(net235),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _2069_ (.A(net235),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _2070_ (.A(net238),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _2071_ (.A(net238),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _2072_ (.A(net236),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _2073_ (.A(net236),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _2074_ (.A(net236),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _2075_ (.A(net236),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _2076_ (.A(net236),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _2077_ (.A(net236),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _2078_ (.A(net238),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _2079_ (.A(net238),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _2080_ (.A(net238),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _2081_ (.A(net239),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _2082_ (.A(net239),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _2083_ (.A(net237),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _2084_ (.A(net237),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _2085_ (.A(net237),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _2086_ (.A(net232),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _2087_ (.A(net232),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _2088_ (.A(net232),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _2089_ (.A(net231),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _2090_ (.A(net233),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _2091_ (.A(net229),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _2092_ (.A(net229),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _2093_ (.A(net229),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _2094_ (.A(net228),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _2095_ (.A(net228),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _2096_ (.A(net228),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _2097_ (.A(net228),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _2098_ (.A(net233),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _2099_ (.A(net231),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _2100_ (.A(net230),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _2101_ (.A(net230),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _2102_ (.A(net230),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _2103_ (.A(net230),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _2104_ (.A(net229),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _2105_ (.A(net232),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _2106_ (.A(net234),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _2107_ (.A(net234),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _2108_ (.A(net226),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _2109_ (.A(net226),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _2110_ (.A(net226),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _2111_ (.A(net227),
    .Y(_0199_));
 sky130_fd_sc_hd__inv_2 _2112_ (.A(net234),
    .Y(_0200_));
 sky130_fd_sc_hd__inv_2 _2113_ (.A(net234),
    .Y(_0201_));
 sky130_fd_sc_hd__inv_2 _2114_ (.A(net236),
    .Y(_0202_));
 sky130_fd_sc_hd__dfrtp_2 _2115_ (.CLK(clknet_leaf_1_clk),
    .D(_0203_),
    .RESET_B(_0000_),
    .Q(\extended_operand[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2116_ (.CLK(clknet_leaf_1_clk),
    .D(_0204_),
    .RESET_B(_0001_),
    .Q(\extended_operand[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2117_ (.CLK(clknet_leaf_1_clk),
    .D(_0205_),
    .RESET_B(_0002_),
    .Q(\extended_operand[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2118_ (.CLK(clknet_leaf_2_clk),
    .D(_0206_),
    .RESET_B(_0003_),
    .Q(\extended_operand[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2119_ (.CLK(clknet_leaf_3_clk),
    .D(_0207_),
    .RESET_B(_0004_),
    .Q(\extended_operand[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2120_ (.CLK(clknet_leaf_3_clk),
    .D(_0208_),
    .RESET_B(_0005_),
    .Q(\extended_operand[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2121_ (.CLK(clknet_leaf_3_clk),
    .D(_0209_),
    .RESET_B(_0006_),
    .Q(\extended_operand[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2122_ (.CLK(clknet_leaf_3_clk),
    .D(_0210_),
    .RESET_B(_0007_),
    .Q(\extended_operand[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2123_ (.CLK(clknet_leaf_3_clk),
    .D(_0211_),
    .RESET_B(_0008_),
    .Q(\extended_operand[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2124_ (.CLK(clknet_leaf_3_clk),
    .D(_0212_),
    .RESET_B(_0009_),
    .Q(\extended_operand[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2125_ (.CLK(clknet_leaf_0_clk),
    .D(_0213_),
    .RESET_B(_0010_),
    .Q(\extended_operand[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2126_ (.CLK(clknet_leaf_0_clk),
    .D(_0214_),
    .RESET_B(_0011_),
    .Q(\extended_operand[11] ));
 sky130_fd_sc_hd__dfrtp_4 _2127_ (.CLK(clknet_leaf_0_clk),
    .D(_0215_),
    .RESET_B(_0012_),
    .Q(\extended_operand[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2128_ (.CLK(clknet_leaf_0_clk),
    .D(_0216_),
    .RESET_B(_0013_),
    .Q(\extended_operand[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2129_ (.CLK(clknet_leaf_23_clk),
    .D(_0217_),
    .RESET_B(_0014_),
    .Q(\extended_operand[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2130_ (.CLK(clknet_leaf_23_clk),
    .D(_0218_),
    .RESET_B(_0015_),
    .Q(\extended_operand[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2131_ (.CLK(clknet_leaf_22_clk),
    .D(_0219_),
    .RESET_B(_0016_),
    .Q(\extended_operand[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2132_ (.CLK(clknet_leaf_22_clk),
    .D(_0220_),
    .RESET_B(_0017_),
    .Q(\extended_operand[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2133_ (.CLK(clknet_leaf_22_clk),
    .D(_0221_),
    .RESET_B(_0018_),
    .Q(\extended_operand[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2134_ (.CLK(clknet_leaf_22_clk),
    .D(_0222_),
    .RESET_B(_0019_),
    .Q(\extended_operand[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2135_ (.CLK(clknet_leaf_21_clk),
    .D(_0223_),
    .RESET_B(_0020_),
    .Q(\extended_operand[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2136_ (.CLK(clknet_leaf_21_clk),
    .D(_0224_),
    .RESET_B(_0021_),
    .Q(\extended_operand[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2137_ (.CLK(clknet_leaf_21_clk),
    .D(_0225_),
    .RESET_B(_0022_),
    .Q(\extended_operand[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2138_ (.CLK(clknet_leaf_21_clk),
    .D(_0226_),
    .RESET_B(_0023_),
    .Q(\extended_operand[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2139_ (.CLK(clknet_leaf_19_clk),
    .D(_0227_),
    .RESET_B(_0024_),
    .Q(\extended_operand[24] ));
 sky130_fd_sc_hd__dfrtp_1 _2140_ (.CLK(clknet_leaf_19_clk),
    .D(_0228_),
    .RESET_B(_0025_),
    .Q(\extended_operand[25] ));
 sky130_fd_sc_hd__dfrtp_1 _2141_ (.CLK(clknet_leaf_19_clk),
    .D(_0229_),
    .RESET_B(_0026_),
    .Q(\extended_operand[26] ));
 sky130_fd_sc_hd__dfrtp_1 _2142_ (.CLK(clknet_leaf_19_clk),
    .D(_0230_),
    .RESET_B(_0027_),
    .Q(\extended_operand[27] ));
 sky130_fd_sc_hd__dfrtp_1 _2143_ (.CLK(clknet_leaf_19_clk),
    .D(_0231_),
    .RESET_B(_0028_),
    .Q(\extended_operand[28] ));
 sky130_fd_sc_hd__dfrtp_1 _2144_ (.CLK(clknet_leaf_19_clk),
    .D(_0232_),
    .RESET_B(_0029_),
    .Q(\extended_operand[29] ));
 sky130_fd_sc_hd__dfrtp_1 _2145_ (.CLK(clknet_leaf_18_clk),
    .D(_0233_),
    .RESET_B(_0030_),
    .Q(\extended_operand[30] ));
 sky130_fd_sc_hd__dfrtp_1 _2146_ (.CLK(clknet_leaf_18_clk),
    .D(_0234_),
    .RESET_B(_0031_),
    .Q(\extended_operand[31] ));
 sky130_fd_sc_hd__dfrtp_1 _2147_ (.CLK(clknet_leaf_14_clk),
    .D(_0235_),
    .RESET_B(_0032_),
    .Q(\partial_sum[63] ));
 sky130_fd_sc_hd__dfrtp_1 _2148_ (.CLK(clknet_leaf_6_clk),
    .D(_0236_),
    .RESET_B(_0033_),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _2149_ (.CLK(clknet_leaf_6_clk),
    .D(_0237_),
    .RESET_B(_0034_),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _2150_ (.CLK(clknet_leaf_9_clk),
    .D(_0238_),
    .RESET_B(_0035_),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_1 _2151_ (.CLK(clknet_leaf_10_clk),
    .D(_0239_),
    .RESET_B(_0036_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _2152_ (.CLK(clknet_leaf_11_clk),
    .D(_0240_),
    .RESET_B(_0037_),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_1 _2153_ (.CLK(clknet_leaf_11_clk),
    .D(_0241_),
    .RESET_B(_0038_),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_1 _2154_ (.CLK(clknet_leaf_12_clk),
    .D(_0242_),
    .RESET_B(_0039_),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_1 _2155_ (.CLK(clknet_leaf_12_clk),
    .D(_0243_),
    .RESET_B(_0040_),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_1 _2156_ (.CLK(clknet_leaf_11_clk),
    .D(_0244_),
    .RESET_B(_0041_),
    .Q(net130));
 sky130_fd_sc_hd__dfrtp_1 _2157_ (.CLK(clknet_leaf_11_clk),
    .D(_0245_),
    .RESET_B(_0042_),
    .Q(net131));
 sky130_fd_sc_hd__dfrtp_1 _2158_ (.CLK(clknet_leaf_10_clk),
    .D(_0246_),
    .RESET_B(_0043_),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _2159_ (.CLK(clknet_leaf_10_clk),
    .D(_0247_),
    .RESET_B(_0044_),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _2160_ (.CLK(clknet_leaf_10_clk),
    .D(_0248_),
    .RESET_B(_0045_),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _2161_ (.CLK(clknet_leaf_6_clk),
    .D(_0249_),
    .RESET_B(_0046_),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _2162_ (.CLK(clknet_leaf_6_clk),
    .D(_0250_),
    .RESET_B(_0047_),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _2163_ (.CLK(clknet_leaf_6_clk),
    .D(_0251_),
    .RESET_B(_0048_),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _2164_ (.CLK(clknet_leaf_5_clk),
    .D(_0252_),
    .RESET_B(_0049_),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _2165_ (.CLK(clknet_leaf_4_clk),
    .D(_0253_),
    .RESET_B(_0050_),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _2166_ (.CLK(clknet_leaf_4_clk),
    .D(_0254_),
    .RESET_B(_0051_),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _2167_ (.CLK(clknet_leaf_4_clk),
    .D(_0255_),
    .RESET_B(_0052_),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _2168_ (.CLK(clknet_leaf_4_clk),
    .D(_0256_),
    .RESET_B(_0053_),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _2169_ (.CLK(clknet_leaf_4_clk),
    .D(_0257_),
    .RESET_B(_0054_),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _2170_ (.CLK(clknet_leaf_4_clk),
    .D(_0258_),
    .RESET_B(_0055_),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _2171_ (.CLK(clknet_leaf_4_clk),
    .D(_0259_),
    .RESET_B(_0056_),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _2172_ (.CLK(clknet_leaf_4_clk),
    .D(_0260_),
    .RESET_B(_0057_),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _2173_ (.CLK(clknet_leaf_4_clk),
    .D(_0261_),
    .RESET_B(_0058_),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _2174_ (.CLK(clknet_leaf_5_clk),
    .D(_0262_),
    .RESET_B(_0059_),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _2175_ (.CLK(clknet_leaf_5_clk),
    .D(_0263_),
    .RESET_B(_0060_),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _2176_ (.CLK(clknet_leaf_5_clk),
    .D(_0264_),
    .RESET_B(_0061_),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _2177_ (.CLK(clknet_leaf_6_clk),
    .D(_0265_),
    .RESET_B(_0062_),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _2178_ (.CLK(clknet_leaf_6_clk),
    .D(_0266_),
    .RESET_B(_0063_),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _2179_ (.CLK(clknet_leaf_6_clk),
    .D(_0267_),
    .RESET_B(_0064_),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _2180_ (.CLK(clknet_leaf_3_clk),
    .D(_0268_),
    .RESET_B(_0065_),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _2181_ (.CLK(clknet_leaf_13_clk),
    .D(_0269_),
    .RESET_B(_0066_),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _2182_ (.CLK(clknet_leaf_17_clk),
    .D(_0270_),
    .RESET_B(_0067_),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _2183_ (.CLK(clknet_leaf_3_clk),
    .D(_0271_),
    .RESET_B(_0068_),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _2184_ (.CLK(clknet_leaf_3_clk),
    .D(_0272_),
    .RESET_B(_0069_),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _2185_ (.CLK(clknet_leaf_3_clk),
    .D(_0273_),
    .RESET_B(_0070_),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _2186_ (.CLK(clknet_leaf_5_clk),
    .D(_0274_),
    .RESET_B(_0071_),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_1 _2187_ (.CLK(clknet_leaf_4_clk),
    .D(_0275_),
    .RESET_B(_0072_),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _2188_ (.CLK(clknet_leaf_3_clk),
    .D(_0276_),
    .RESET_B(_0073_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _2189_ (.CLK(clknet_leaf_3_clk),
    .D(_0277_),
    .RESET_B(_0074_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _2190_ (.CLK(clknet_leaf_0_clk),
    .D(_0278_),
    .RESET_B(_0075_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _2191_ (.CLK(clknet_leaf_0_clk),
    .D(_0279_),
    .RESET_B(_0076_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_1 _2192_ (.CLK(clknet_leaf_20_clk),
    .D(_0280_),
    .RESET_B(_0077_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_1 _2193_ (.CLK(clknet_leaf_0_clk),
    .D(_0281_),
    .RESET_B(_0078_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_1 _2194_ (.CLK(clknet_leaf_0_clk),
    .D(_0282_),
    .RESET_B(_0079_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_1 _2195_ (.CLK(clknet_leaf_22_clk),
    .D(_0283_),
    .RESET_B(_0080_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_1 _2196_ (.CLK(clknet_leaf_23_clk),
    .D(_0284_),
    .RESET_B(_0081_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_1 _2197_ (.CLK(clknet_leaf_22_clk),
    .D(_0285_),
    .RESET_B(_0082_),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_1 _2198_ (.CLK(clknet_leaf_22_clk),
    .D(_0286_),
    .RESET_B(_0083_),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_1 _2199_ (.CLK(clknet_leaf_21_clk),
    .D(_0287_),
    .RESET_B(_0084_),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_1 _2200_ (.CLK(clknet_leaf_21_clk),
    .D(_0288_),
    .RESET_B(_0085_),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_1 _2201_ (.CLK(clknet_leaf_21_clk),
    .D(_0289_),
    .RESET_B(_0086_),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_1 _2202_ (.CLK(clknet_leaf_21_clk),
    .D(_0290_),
    .RESET_B(_0087_),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_1 _2203_ (.CLK(clknet_leaf_17_clk),
    .D(_0291_),
    .RESET_B(_0088_),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_1 _2204_ (.CLK(clknet_leaf_17_clk),
    .D(_0292_),
    .RESET_B(_0089_),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_1 _2205_ (.CLK(clknet_leaf_17_clk),
    .D(_0293_),
    .RESET_B(_0090_),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_1 _2206_ (.CLK(clknet_leaf_17_clk),
    .D(_0294_),
    .RESET_B(_0091_),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_1 _2207_ (.CLK(clknet_leaf_17_clk),
    .D(_0295_),
    .RESET_B(_0092_),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_1 _2208_ (.CLK(clknet_leaf_17_clk),
    .D(_0296_),
    .RESET_B(_0093_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_1 _2209_ (.CLK(clknet_leaf_17_clk),
    .D(_0297_),
    .RESET_B(_0094_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_1 _2210_ (.CLK(clknet_leaf_18_clk),
    .D(_0298_),
    .RESET_B(_0095_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_1 _2211_ (.CLK(clknet_leaf_18_clk),
    .D(_0299_),
    .RESET_B(_0096_),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_1 _2212_ (.CLK(clknet_leaf_3_clk),
    .D(_0300_),
    .RESET_B(_0097_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _2213_ (.CLK(clknet_leaf_2_clk),
    .D(_0301_),
    .RESET_B(_0098_),
    .Q(\partial_sum[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2214_ (.CLK(clknet_leaf_2_clk),
    .D(_0302_),
    .RESET_B(_0099_),
    .Q(\partial_sum[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2215_ (.CLK(clknet_leaf_2_clk),
    .D(_0303_),
    .RESET_B(_0100_),
    .Q(\partial_sum[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2216_ (.CLK(clknet_leaf_2_clk),
    .D(_0304_),
    .RESET_B(_0101_),
    .Q(\partial_sum[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2217_ (.CLK(clknet_leaf_2_clk),
    .D(_0305_),
    .RESET_B(_0102_),
    .Q(\partial_sum[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2218_ (.CLK(clknet_leaf_7_clk),
    .D(_0306_),
    .RESET_B(_0103_),
    .Q(\partial_sum[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2219_ (.CLK(clknet_leaf_7_clk),
    .D(_0307_),
    .RESET_B(_0104_),
    .Q(\partial_sum[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2220_ (.CLK(clknet_leaf_5_clk),
    .D(_0308_),
    .RESET_B(_0105_),
    .Q(\partial_sum[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2221_ (.CLK(clknet_leaf_2_clk),
    .D(_0309_),
    .RESET_B(_0106_),
    .Q(\partial_sum[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2222_ (.CLK(clknet_leaf_1_clk),
    .D(_0310_),
    .RESET_B(_0107_),
    .Q(\partial_sum[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2223_ (.CLK(clknet_leaf_1_clk),
    .D(_0311_),
    .RESET_B(_0108_),
    .Q(\partial_sum[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2224_ (.CLK(clknet_leaf_1_clk),
    .D(_0312_),
    .RESET_B(_0109_),
    .Q(\partial_sum[11] ));
 sky130_fd_sc_hd__dfrtp_2 _2225_ (.CLK(clknet_leaf_1_clk),
    .D(_0313_),
    .RESET_B(_0110_),
    .Q(\partial_sum[12] ));
 sky130_fd_sc_hd__dfrtp_2 _2226_ (.CLK(clknet_leaf_1_clk),
    .D(_0314_),
    .RESET_B(_0111_),
    .Q(\partial_sum[13] ));
 sky130_fd_sc_hd__dfrtp_2 _2227_ (.CLK(clknet_leaf_1_clk),
    .D(_0315_),
    .RESET_B(_0112_),
    .Q(\partial_sum[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2228_ (.CLK(clknet_leaf_23_clk),
    .D(_0316_),
    .RESET_B(_0113_),
    .Q(\partial_sum[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2229_ (.CLK(clknet_leaf_23_clk),
    .D(_0317_),
    .RESET_B(_0114_),
    .Q(\partial_sum[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2230_ (.CLK(clknet_leaf_22_clk),
    .D(_0318_),
    .RESET_B(_0115_),
    .Q(\partial_sum[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2231_ (.CLK(clknet_leaf_22_clk),
    .D(_0319_),
    .RESET_B(_0116_),
    .Q(\partial_sum[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2232_ (.CLK(clknet_leaf_21_clk),
    .D(_0320_),
    .RESET_B(_0117_),
    .Q(\partial_sum[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2233_ (.CLK(clknet_leaf_21_clk),
    .D(_0321_),
    .RESET_B(_0118_),
    .Q(\partial_sum[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2234_ (.CLK(clknet_leaf_20_clk),
    .D(_0322_),
    .RESET_B(_0119_),
    .Q(\partial_sum[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2235_ (.CLK(clknet_leaf_20_clk),
    .D(_0323_),
    .RESET_B(_0120_),
    .Q(\partial_sum[22] ));
 sky130_fd_sc_hd__dfrtp_2 _2236_ (.CLK(clknet_leaf_20_clk),
    .D(_0324_),
    .RESET_B(_0121_),
    .Q(\partial_sum[23] ));
 sky130_fd_sc_hd__dfrtp_4 _2237_ (.CLK(clknet_leaf_19_clk),
    .D(_0325_),
    .RESET_B(_0122_),
    .Q(\partial_sum[24] ));
 sky130_fd_sc_hd__dfrtp_4 _2238_ (.CLK(clknet_leaf_20_clk),
    .D(_0326_),
    .RESET_B(_0123_),
    .Q(\partial_sum[25] ));
 sky130_fd_sc_hd__dfrtp_4 _2239_ (.CLK(clknet_leaf_16_clk),
    .D(_0327_),
    .RESET_B(_0124_),
    .Q(\partial_sum[26] ));
 sky130_fd_sc_hd__dfrtp_2 _2240_ (.CLK(clknet_leaf_16_clk),
    .D(_0328_),
    .RESET_B(_0125_),
    .Q(\partial_sum[27] ));
 sky130_fd_sc_hd__dfrtp_2 _2241_ (.CLK(clknet_leaf_18_clk),
    .D(_0329_),
    .RESET_B(_0126_),
    .Q(\partial_sum[28] ));
 sky130_fd_sc_hd__dfrtp_2 _2242_ (.CLK(clknet_leaf_18_clk),
    .D(_0330_),
    .RESET_B(_0127_),
    .Q(\partial_sum[29] ));
 sky130_fd_sc_hd__dfrtp_2 _2243_ (.CLK(clknet_leaf_18_clk),
    .D(_0331_),
    .RESET_B(_0128_),
    .Q(\partial_sum[30] ));
 sky130_fd_sc_hd__dfrtp_2 _2244_ (.CLK(clknet_leaf_18_clk),
    .D(_0332_),
    .RESET_B(_0129_),
    .Q(\partial_sum[31] ));
 sky130_fd_sc_hd__dfrtp_2 _2245_ (.CLK(clknet_leaf_18_clk),
    .D(_0333_),
    .RESET_B(_0130_),
    .Q(\partial_sum[32] ));
 sky130_fd_sc_hd__dfrtp_1 _2246_ (.CLK(clknet_leaf_17_clk),
    .D(_0334_),
    .RESET_B(_0131_),
    .Q(\partial_sum[33] ));
 sky130_fd_sc_hd__dfrtp_1 _2247_ (.CLK(clknet_leaf_17_clk),
    .D(_0335_),
    .RESET_B(_0132_),
    .Q(\partial_sum[34] ));
 sky130_fd_sc_hd__dfrtp_1 _2248_ (.CLK(clknet_leaf_16_clk),
    .D(_0336_),
    .RESET_B(_0133_),
    .Q(\partial_sum[35] ));
 sky130_fd_sc_hd__dfrtp_1 _2249_ (.CLK(clknet_leaf_16_clk),
    .D(_0337_),
    .RESET_B(_0134_),
    .Q(\partial_sum[36] ));
 sky130_fd_sc_hd__dfrtp_1 _2250_ (.CLK(clknet_leaf_16_clk),
    .D(_0338_),
    .RESET_B(_0135_),
    .Q(\partial_sum[37] ));
 sky130_fd_sc_hd__dfrtp_1 _2251_ (.CLK(clknet_leaf_15_clk),
    .D(_0339_),
    .RESET_B(_0136_),
    .Q(\partial_sum[38] ));
 sky130_fd_sc_hd__dfrtp_1 _2252_ (.CLK(clknet_leaf_20_clk),
    .D(_0340_),
    .RESET_B(_0137_),
    .Q(\partial_sum[39] ));
 sky130_fd_sc_hd__dfrtp_1 _2253_ (.CLK(clknet_leaf_20_clk),
    .D(_0341_),
    .RESET_B(_0138_),
    .Q(\partial_sum[40] ));
 sky130_fd_sc_hd__dfrtp_1 _2254_ (.CLK(clknet_leaf_20_clk),
    .D(_0342_),
    .RESET_B(_0139_),
    .Q(\partial_sum[41] ));
 sky130_fd_sc_hd__dfrtp_1 _2255_ (.CLK(clknet_leaf_20_clk),
    .D(_0343_),
    .RESET_B(_0140_),
    .Q(\partial_sum[42] ));
 sky130_fd_sc_hd__dfrtp_1 _2256_ (.CLK(clknet_leaf_1_clk),
    .D(_0344_),
    .RESET_B(_0141_),
    .Q(\partial_sum[43] ));
 sky130_fd_sc_hd__dfrtp_1 _2257_ (.CLK(clknet_leaf_20_clk),
    .D(_0345_),
    .RESET_B(_0142_),
    .Q(\partial_sum[44] ));
 sky130_fd_sc_hd__dfrtp_1 _2258_ (.CLK(clknet_leaf_20_clk),
    .D(_0346_),
    .RESET_B(_0143_),
    .Q(\partial_sum[45] ));
 sky130_fd_sc_hd__dfrtp_1 _2259_ (.CLK(clknet_leaf_15_clk),
    .D(_0347_),
    .RESET_B(_0144_),
    .Q(\partial_sum[46] ));
 sky130_fd_sc_hd__dfrtp_1 _2260_ (.CLK(clknet_leaf_15_clk),
    .D(_0348_),
    .RESET_B(_0145_),
    .Q(\partial_sum[47] ));
 sky130_fd_sc_hd__dfrtp_1 _2261_ (.CLK(clknet_leaf_14_clk),
    .D(_0349_),
    .RESET_B(_0146_),
    .Q(\partial_sum[48] ));
 sky130_fd_sc_hd__dfrtp_1 _2262_ (.CLK(clknet_leaf_14_clk),
    .D(_0350_),
    .RESET_B(_0147_),
    .Q(\partial_sum[49] ));
 sky130_fd_sc_hd__dfrtp_1 _2263_ (.CLK(clknet_leaf_8_clk),
    .D(_0351_),
    .RESET_B(_0148_),
    .Q(\partial_sum[50] ));
 sky130_fd_sc_hd__dfrtp_1 _2264_ (.CLK(clknet_leaf_14_clk),
    .D(_0352_),
    .RESET_B(_0149_),
    .Q(\partial_sum[51] ));
 sky130_fd_sc_hd__dfrtp_2 _2265_ (.CLK(clknet_leaf_14_clk),
    .D(_0353_),
    .RESET_B(_0150_),
    .Q(\partial_sum[52] ));
 sky130_fd_sc_hd__dfrtp_1 _2266_ (.CLK(clknet_leaf_17_clk),
    .D(_0354_),
    .RESET_B(_0151_),
    .Q(\partial_sum[53] ));
 sky130_fd_sc_hd__dfrtp_1 _2267_ (.CLK(clknet_leaf_13_clk),
    .D(_0355_),
    .RESET_B(_0152_),
    .Q(\partial_sum[54] ));
 sky130_fd_sc_hd__dfrtp_1 _2268_ (.CLK(clknet_leaf_13_clk),
    .D(_0356_),
    .RESET_B(_0153_),
    .Q(\partial_sum[55] ));
 sky130_fd_sc_hd__dfrtp_2 _2269_ (.CLK(clknet_leaf_13_clk),
    .D(_0357_),
    .RESET_B(_0154_),
    .Q(\partial_sum[56] ));
 sky130_fd_sc_hd__dfrtp_2 _2270_ (.CLK(clknet_leaf_13_clk),
    .D(_0358_),
    .RESET_B(_0155_),
    .Q(\partial_sum[57] ));
 sky130_fd_sc_hd__dfrtp_1 _2271_ (.CLK(clknet_leaf_12_clk),
    .D(_0359_),
    .RESET_B(_0156_),
    .Q(\partial_sum[58] ));
 sky130_fd_sc_hd__dfrtp_1 _2272_ (.CLK(clknet_leaf_12_clk),
    .D(_0360_),
    .RESET_B(_0157_),
    .Q(\partial_sum[59] ));
 sky130_fd_sc_hd__dfrtp_1 _2273_ (.CLK(clknet_leaf_12_clk),
    .D(_0361_),
    .RESET_B(_0158_),
    .Q(\partial_sum[60] ));
 sky130_fd_sc_hd__dfrtp_1 _2274_ (.CLK(clknet_leaf_11_clk),
    .D(_0362_),
    .RESET_B(_0159_),
    .Q(\partial_sum[61] ));
 sky130_fd_sc_hd__dfrtp_1 _2275_ (.CLK(clknet_leaf_9_clk),
    .D(_0363_),
    .RESET_B(_0160_),
    .Q(\partial_sum[62] ));
 sky130_fd_sc_hd__dfrtp_2 _2276_ (.CLK(clknet_leaf_9_clk),
    .D(_0364_),
    .RESET_B(_0161_),
    .Q(\current_multiplier[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2277_ (.CLK(clknet_leaf_10_clk),
    .D(_0365_),
    .RESET_B(_0162_),
    .Q(\current_multiplier[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2278_ (.CLK(clknet_leaf_10_clk),
    .D(_0366_),
    .RESET_B(_0163_),
    .Q(\current_multiplier[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2279_ (.CLK(clknet_leaf_10_clk),
    .D(_0367_),
    .RESET_B(_0164_),
    .Q(\current_multiplier[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2280_ (.CLK(clknet_leaf_10_clk),
    .D(_0368_),
    .RESET_B(_0165_),
    .Q(\current_multiplier[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2281_ (.CLK(clknet_leaf_11_clk),
    .D(_0369_),
    .RESET_B(_0166_),
    .Q(\current_multiplier[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2282_ (.CLK(clknet_leaf_11_clk),
    .D(_0370_),
    .RESET_B(_0167_),
    .Q(\current_multiplier[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2283_ (.CLK(clknet_leaf_11_clk),
    .D(_0371_),
    .RESET_B(_0168_),
    .Q(\current_multiplier[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2284_ (.CLK(clknet_leaf_11_clk),
    .D(_0372_),
    .RESET_B(_0169_),
    .Q(\current_multiplier[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2285_ (.CLK(clknet_leaf_11_clk),
    .D(_0373_),
    .RESET_B(_0170_),
    .Q(\current_multiplier[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2286_ (.CLK(clknet_leaf_10_clk),
    .D(_0374_),
    .RESET_B(_0171_),
    .Q(\current_multiplier[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2287_ (.CLK(clknet_leaf_10_clk),
    .D(_0375_),
    .RESET_B(_0172_),
    .Q(\current_multiplier[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2288_ (.CLK(clknet_leaf_10_clk),
    .D(_0376_),
    .RESET_B(_0173_),
    .Q(\current_multiplier[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2289_ (.CLK(clknet_leaf_6_clk),
    .D(_0377_),
    .RESET_B(_0174_),
    .Q(\current_multiplier[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2290_ (.CLK(clknet_leaf_9_clk),
    .D(_0378_),
    .RESET_B(_0175_),
    .Q(\current_multiplier[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2291_ (.CLK(clknet_leaf_5_clk),
    .D(_0379_),
    .RESET_B(_0176_),
    .Q(\current_multiplier[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2292_ (.CLK(clknet_leaf_5_clk),
    .D(_0380_),
    .RESET_B(_0177_),
    .Q(\current_multiplier[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2293_ (.CLK(clknet_leaf_4_clk),
    .D(_0381_),
    .RESET_B(_0178_),
    .Q(\current_multiplier[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2294_ (.CLK(clknet_leaf_4_clk),
    .D(_0382_),
    .RESET_B(_0179_),
    .Q(\current_multiplier[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2295_ (.CLK(clknet_leaf_4_clk),
    .D(_0383_),
    .RESET_B(_0180_),
    .Q(\current_multiplier[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2296_ (.CLK(clknet_leaf_4_clk),
    .D(_0384_),
    .RESET_B(_0181_),
    .Q(\current_multiplier[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2297_ (.CLK(clknet_leaf_4_clk),
    .D(_0385_),
    .RESET_B(_0182_),
    .Q(\current_multiplier[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2298_ (.CLK(clknet_leaf_4_clk),
    .D(_0386_),
    .RESET_B(_0183_),
    .Q(\current_multiplier[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2299_ (.CLK(clknet_leaf_4_clk),
    .D(_0387_),
    .RESET_B(_0184_),
    .Q(\current_multiplier[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2300_ (.CLK(clknet_leaf_4_clk),
    .D(_0388_),
    .RESET_B(_0185_),
    .Q(\current_multiplier[24] ));
 sky130_fd_sc_hd__dfrtp_1 _2301_ (.CLK(clknet_leaf_4_clk),
    .D(_0389_),
    .RESET_B(_0186_),
    .Q(\current_multiplier[25] ));
 sky130_fd_sc_hd__dfrtp_1 _2302_ (.CLK(clknet_leaf_5_clk),
    .D(_0390_),
    .RESET_B(_0187_),
    .Q(\current_multiplier[26] ));
 sky130_fd_sc_hd__dfrtp_1 _2303_ (.CLK(clknet_leaf_5_clk),
    .D(_0391_),
    .RESET_B(_0188_),
    .Q(\current_multiplier[27] ));
 sky130_fd_sc_hd__dfrtp_1 _2304_ (.CLK(clknet_leaf_6_clk),
    .D(_0392_),
    .RESET_B(_0189_),
    .Q(\current_multiplier[28] ));
 sky130_fd_sc_hd__dfrtp_1 _2305_ (.CLK(clknet_leaf_6_clk),
    .D(_0393_),
    .RESET_B(_0190_),
    .Q(\current_multiplier[29] ));
 sky130_fd_sc_hd__dfrtp_1 _2306_ (.CLK(clknet_leaf_6_clk),
    .D(_0394_),
    .RESET_B(_0191_),
    .Q(\current_multiplier[30] ));
 sky130_fd_sc_hd__dfrtp_1 _2307_ (.CLK(clknet_leaf_4_clk),
    .D(_0395_),
    .RESET_B(_0192_),
    .Q(\current_multiplier[31] ));
 sky130_fd_sc_hd__dfrtp_1 _2308_ (.CLK(clknet_leaf_6_clk),
    .D(_0396_),
    .RESET_B(_0193_),
    .Q(last_bit));
 sky130_fd_sc_hd__dfrtp_1 _2309_ (.CLK(clknet_leaf_8_clk),
    .D(_0397_),
    .RESET_B(_0194_),
    .Q(\iteration_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2310_ (.CLK(clknet_leaf_8_clk),
    .D(_0398_),
    .RESET_B(_0195_),
    .Q(\iteration_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2311_ (.CLK(clknet_leaf_8_clk),
    .D(_0399_),
    .RESET_B(_0196_),
    .Q(\iteration_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2312_ (.CLK(clknet_leaf_8_clk),
    .D(_0400_),
    .RESET_B(_0197_),
    .Q(\iteration_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2313_ (.CLK(clknet_leaf_7_clk),
    .D(_0401_),
    .RESET_B(_0198_),
    .Q(\iteration_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2314_ (.CLK(clknet_leaf_7_clk),
    .D(_0402_),
    .RESET_B(_0199_),
    .Q(\iteration_count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2315_ (.CLK(clknet_leaf_8_clk),
    .D(\next_state[0] ),
    .RESET_B(_0200_),
    .Q(\current_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2316_ (.CLK(clknet_leaf_9_clk),
    .D(\next_state[1] ),
    .RESET_B(_0201_),
    .Q(\current_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2317_ (.CLK(clknet_leaf_9_clk),
    .D(\next_state[2] ),
    .RESET_B(_0202_),
    .Q(\current_state[2] ));
 sky130_fd_sc_hd__buf_1 input1 (.A(M[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(M[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(M[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(M[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(M[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(M[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(M[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(M[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(M[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(M[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(M[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(M[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(M[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(M[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(M[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(M[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(M[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(M[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(M[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(M[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(M[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(M[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(M[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(M[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(M[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(M[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(M[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(M[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(M[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(M[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(M[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(M[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(Q[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(Q[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(Q[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(Q[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(Q[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(Q[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(Q[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(Q[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(Q[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(Q[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(Q[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(Q[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(Q[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(Q[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(Q[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(Q[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(Q[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(Q[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(Q[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(Q[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(Q[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(Q[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(Q[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(Q[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(Q[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(Q[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(Q[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(Q[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(Q[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(Q[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(Q[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(Q[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(rst),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(start),
    .X(net66));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(done));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(result[0]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(result[10]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(result[11]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(result[12]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(result[13]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(result[14]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(result[15]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(result[16]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(result[17]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(result[18]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(result[19]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(result[1]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(result[20]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(result[21]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(result[22]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(result[23]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(result[24]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(result[25]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(result[26]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(result[27]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(result[28]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(result[29]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(result[2]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(result[30]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(result[31]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(result[32]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(result[33]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(result[34]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(result[35]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(result[36]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(result[37]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(result[38]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(result[39]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(result[3]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(result[40]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(result[41]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(result[42]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(result[43]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(result[44]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(result[45]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(result[46]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(result[47]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(result[48]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(result[49]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(result[4]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(result[50]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(result[51]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(result[52]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(result[53]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(result[54]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(result[55]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(result[56]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(result[57]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(result[58]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(result[59]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(result[5]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(result[60]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(result[61]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(result[62]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(result[63]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(result[6]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(result[7]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(result[8]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(result[9]));
 sky130_fd_sc_hd__clkbuf_1 wire132 (.A(_0987_),
    .X(net132));
 sky130_fd_sc_hd__buf_2 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_2 fanout134 (.A(_0852_),
    .X(net134));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 fanout136 (.A(net140),
    .X(net136));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(net140),
    .X(net137));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net140),
    .X(net138));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 fanout140 (.A(_0852_),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 fanout141 (.A(_0494_),
    .X(net141));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(net144),
    .X(net142));
 sky130_fd_sc_hd__buf_2 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(_0493_),
    .X(net144));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_2 fanout146 (.A(_0493_),
    .X(net146));
 sky130_fd_sc_hd__buf_2 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_2 fanout148 (.A(_0493_),
    .X(net148));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(_0837_),
    .X(net149));
 sky130_fd_sc_hd__buf_2 fanout150 (.A(_0792_),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 fanout151 (.A(_0792_),
    .X(net151));
 sky130_fd_sc_hd__buf_2 fanout152 (.A(_0792_),
    .X(net152));
 sky130_fd_sc_hd__buf_1 fanout153 (.A(_0792_),
    .X(net153));
 sky130_fd_sc_hd__buf_2 fanout154 (.A(_0786_),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(_0786_),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(_0786_),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 fanout157 (.A(_0786_),
    .X(net157));
 sky130_fd_sc_hd__buf_2 fanout158 (.A(net161),
    .X(net158));
 sky130_fd_sc_hd__buf_2 fanout159 (.A(net161),
    .X(net159));
 sky130_fd_sc_hd__buf_2 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 fanout161 (.A(_0785_),
    .X(net161));
 sky130_fd_sc_hd__buf_2 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__buf_2 fanout163 (.A(_0785_),
    .X(net163));
 sky130_fd_sc_hd__buf_2 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 fanout165 (.A(_0785_),
    .X(net165));
 sky130_fd_sc_hd__buf_2 fanout166 (.A(net171),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 fanout167 (.A(net170),
    .X(net167));
 sky130_fd_sc_hd__buf_1 fanout168 (.A(net170),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 fanout171 (.A(_0700_),
    .X(net171));
 sky130_fd_sc_hd__buf_2 fanout172 (.A(net174),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 fanout173 (.A(_0700_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 fanout174 (.A(_0700_),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(net179),
    .X(net175));
 sky130_fd_sc_hd__buf_2 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 fanout177 (.A(net179),
    .X(net177));
 sky130_fd_sc_hd__buf_2 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_2 fanout179 (.A(_0699_),
    .X(net179));
 sky130_fd_sc_hd__buf_2 fanout180 (.A(net182),
    .X(net180));
 sky130_fd_sc_hd__buf_2 fanout181 (.A(_0699_),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 fanout182 (.A(_0699_),
    .X(net182));
 sky130_fd_sc_hd__buf_2 fanout183 (.A(net186),
    .X(net183));
 sky130_fd_sc_hd__buf_2 fanout184 (.A(net186),
    .X(net184));
 sky130_fd_sc_hd__buf_2 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__buf_2 fanout186 (.A(_0849_),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(_0848_),
    .X(net187));
 sky130_fd_sc_hd__buf_2 fanout188 (.A(_0848_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(_0848_),
    .X(net189));
 sky130_fd_sc_hd__buf_2 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(net194),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net194),
    .X(net192));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 fanout194 (.A(_0847_),
    .X(net194));
 sky130_fd_sc_hd__buf_2 fanout195 (.A(net198),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 fanout196 (.A(net198),
    .X(net196));
 sky130_fd_sc_hd__buf_2 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 fanout198 (.A(net211),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 fanout200 (.A(net211),
    .X(net200));
 sky130_fd_sc_hd__buf_2 fanout201 (.A(net207),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 fanout203 (.A(net206),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 fanout207 (.A(net211),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 fanout211 (.A(_0790_),
    .X(net211));
 sky130_fd_sc_hd__buf_2 fanout212 (.A(\current_state[2] ),
    .X(net212));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(net215),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_4 fanout215 (.A(net224),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(net218),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__buf_2 fanout218 (.A(net224),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net224),
    .X(net219));
 sky130_fd_sc_hd__buf_2 fanout220 (.A(net224),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(net223),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net224),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_2 fanout224 (.A(net65),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net227),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__buf_2 fanout227 (.A(net240),
    .X(net227));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__buf_4 fanout229 (.A(net233),
    .X(net229));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(net232),
    .X(net230));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__buf_2 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 fanout233 (.A(net240),
    .X(net233));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(net240),
    .X(net234));
 sky130_fd_sc_hd__buf_2 fanout235 (.A(net240),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(net239),
    .X(net236));
 sky130_fd_sc_hd__buf_2 fanout237 (.A(net239),
    .X(net237));
 sky130_fd_sc_hd__buf_4 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 fanout240 (.A(net65),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload0 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__inv_8 clkload1 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinv_8 clkload2 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__inv_8 clkload4 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__inv_12 clkload6 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__inv_8 clkload7 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__inv_8 clkload8 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkinv_8 clkload9 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__inv_12 clkload10 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload11 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload12 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload13 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_4 clkload14 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinv_4 clkload15 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkinv_4 clkload16 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__inv_6 clkload17 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_4 clkload18 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload19 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__bufinv_16 clkload20 (.A(clknet_leaf_19_clk));
endmodule
