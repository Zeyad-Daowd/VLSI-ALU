module sequential_multiplier_shift_accumulate_route (clk,
    done,
    rst,
    multiplicand,
    multiplier,
    product);
 input clk;
 output done;
 input rst;
 input [31:0] multiplicand;
 input [31:0] multiplier;
 output [63:0] product;

 wire \A[0] ;
 wire \A[10] ;
 wire \A[11] ;
 wire \A[12] ;
 wire \A[13] ;
 wire \A[14] ;
 wire \A[15] ;
 wire \A[16] ;
 wire \A[17] ;
 wire \A[18] ;
 wire \A[19] ;
 wire \A[1] ;
 wire \A[20] ;
 wire \A[21] ;
 wire \A[22] ;
 wire \A[23] ;
 wire \A[24] ;
 wire \A[25] ;
 wire \A[26] ;
 wire \A[27] ;
 wire \A[28] ;
 wire \A[29] ;
 wire \A[2] ;
 wire \A[30] ;
 wire \A[31] ;
 wire \A[32] ;
 wire \A[33] ;
 wire \A[34] ;
 wire \A[35] ;
 wire \A[36] ;
 wire \A[37] ;
 wire \A[38] ;
 wire \A[39] ;
 wire \A[3] ;
 wire \A[40] ;
 wire \A[41] ;
 wire \A[42] ;
 wire \A[43] ;
 wire \A[44] ;
 wire \A[45] ;
 wire \A[46] ;
 wire \A[47] ;
 wire \A[48] ;
 wire \A[49] ;
 wire \A[4] ;
 wire \A[50] ;
 wire \A[51] ;
 wire \A[52] ;
 wire \A[53] ;
 wire \A[54] ;
 wire \A[55] ;
 wire \A[56] ;
 wire \A[57] ;
 wire \A[58] ;
 wire \A[59] ;
 wire \A[5] ;
 wire \A[60] ;
 wire \A[61] ;
 wire \A[62] ;
 wire \A[6] ;
 wire \A[7] ;
 wire \A[8] ;
 wire \A[9] ;
 wire \M[0] ;
 wire \M[10] ;
 wire \M[11] ;
 wire \M[12] ;
 wire \M[13] ;
 wire \M[14] ;
 wire \M[15] ;
 wire \M[16] ;
 wire \M[17] ;
 wire \M[18] ;
 wire \M[19] ;
 wire \M[1] ;
 wire \M[20] ;
 wire \M[21] ;
 wire \M[22] ;
 wire \M[23] ;
 wire \M[24] ;
 wire \M[25] ;
 wire \M[26] ;
 wire \M[27] ;
 wire \M[28] ;
 wire \M[29] ;
 wire \M[2] ;
 wire \M[30] ;
 wire \M[31] ;
 wire \M[3] ;
 wire \M[4] ;
 wire \M[5] ;
 wire \M[6] ;
 wire \M[7] ;
 wire \M[8] ;
 wire \M[9] ;
 wire \Q[0] ;
 wire \Q[10] ;
 wire \Q[11] ;
 wire \Q[12] ;
 wire \Q[13] ;
 wire \Q[14] ;
 wire \Q[15] ;
 wire \Q[16] ;
 wire \Q[17] ;
 wire \Q[18] ;
 wire \Q[19] ;
 wire \Q[1] ;
 wire \Q[20] ;
 wire \Q[21] ;
 wire \Q[22] ;
 wire \Q[23] ;
 wire \Q[24] ;
 wire \Q[25] ;
 wire \Q[26] ;
 wire \Q[27] ;
 wire \Q[28] ;
 wire \Q[29] ;
 wire \Q[2] ;
 wire \Q[30] ;
 wire \Q[31] ;
 wire \Q[3] ;
 wire \Q[4] ;
 wire \Q[5] ;
 wire \Q[6] ;
 wire \Q[7] ;
 wire \Q[8] ;
 wire \Q[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire \abs_multiplicand[0] ;
 wire \abs_multiplicand[10] ;
 wire \abs_multiplicand[11] ;
 wire \abs_multiplicand[12] ;
 wire \abs_multiplicand[13] ;
 wire \abs_multiplicand[14] ;
 wire \abs_multiplicand[15] ;
 wire \abs_multiplicand[16] ;
 wire \abs_multiplicand[17] ;
 wire \abs_multiplicand[18] ;
 wire \abs_multiplicand[19] ;
 wire \abs_multiplicand[1] ;
 wire \abs_multiplicand[20] ;
 wire \abs_multiplicand[21] ;
 wire \abs_multiplicand[22] ;
 wire \abs_multiplicand[23] ;
 wire \abs_multiplicand[24] ;
 wire \abs_multiplicand[25] ;
 wire \abs_multiplicand[26] ;
 wire \abs_multiplicand[27] ;
 wire \abs_multiplicand[28] ;
 wire \abs_multiplicand[29] ;
 wire \abs_multiplicand[2] ;
 wire \abs_multiplicand[30] ;
 wire \abs_multiplicand[31] ;
 wire \abs_multiplicand[3] ;
 wire \abs_multiplicand[4] ;
 wire \abs_multiplicand[5] ;
 wire \abs_multiplicand[6] ;
 wire \abs_multiplicand[7] ;
 wire \abs_multiplicand[8] ;
 wire \abs_multiplicand[9] ;
 wire \abs_multiplier[0] ;
 wire \abs_multiplier[10] ;
 wire \abs_multiplier[11] ;
 wire \abs_multiplier[12] ;
 wire \abs_multiplier[13] ;
 wire \abs_multiplier[14] ;
 wire \abs_multiplier[15] ;
 wire \abs_multiplier[16] ;
 wire \abs_multiplier[17] ;
 wire \abs_multiplier[18] ;
 wire \abs_multiplier[19] ;
 wire \abs_multiplier[1] ;
 wire \abs_multiplier[20] ;
 wire \abs_multiplier[21] ;
 wire \abs_multiplier[22] ;
 wire \abs_multiplier[23] ;
 wire \abs_multiplier[24] ;
 wire \abs_multiplier[25] ;
 wire \abs_multiplier[26] ;
 wire \abs_multiplier[27] ;
 wire \abs_multiplier[28] ;
 wire \abs_multiplier[29] ;
 wire \abs_multiplier[2] ;
 wire \abs_multiplier[30] ;
 wire \abs_multiplier[31] ;
 wire \abs_multiplier[3] ;
 wire \abs_multiplier[4] ;
 wire \abs_multiplier[5] ;
 wire \abs_multiplier[6] ;
 wire \abs_multiplier[7] ;
 wire \abs_multiplier[8] ;
 wire \abs_multiplier[9] ;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \count[4] ;
 wire \count[5] ;
 wire sign;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;

 sky130_fd_sc_hd__inv_2 _1152_ (.A(\A[61] ),
    .Y(_0870_));
 sky130_fd_sc_hd__inv_2 _1153_ (.A(\A[54] ),
    .Y(_0871_));
 sky130_fd_sc_hd__inv_2 _1154_ (.A(\A[1] ),
    .Y(_0872_));
 sky130_fd_sc_hd__clkinv_16 _1155_ (.A(\count[5] ),
    .Y(_0873_));
 sky130_fd_sc_hd__inv_2 _1156_ (.A(net26),
    .Y(_0874_));
 sky130_fd_sc_hd__inv_2 _1157_ (.A(net117),
    .Y(_0875_));
 sky130_fd_sc_hd__inv_2 _1158_ (.A(net99),
    .Y(_0876_));
 sky130_fd_sc_hd__inv_2 _1159_ (.A(\Q[28] ),
    .Y(_0877_));
 sky130_fd_sc_hd__inv_2 _1160_ (.A(\Q[24] ),
    .Y(_0878_));
 sky130_fd_sc_hd__inv_2 _1161_ (.A(\Q[22] ),
    .Y(_0879_));
 sky130_fd_sc_hd__inv_2 _1162_ (.A(\Q[13] ),
    .Y(_0880_));
 sky130_fd_sc_hd__inv_2 _1163_ (.A(\Q[10] ),
    .Y(_0881_));
 sky130_fd_sc_hd__inv_2 _1164_ (.A(\Q[4] ),
    .Y(_0882_));
 sky130_fd_sc_hd__inv_2 _1165_ (.A(\M[1] ),
    .Y(_0883_));
 sky130_fd_sc_hd__inv_2 _1166_ (.A(net9),
    .Y(_0884_));
 sky130_fd_sc_hd__inv_2 _1167_ (.A(net22),
    .Y(_0885_));
 sky130_fd_sc_hd__inv_2 _1168_ (.A(net41),
    .Y(_0886_));
 sky130_fd_sc_hd__inv_2 _1169_ (.A(net50),
    .Y(_0887_));
 sky130_fd_sc_hd__inv_2 _1170_ (.A(\abs_multiplicand[31] ),
    .Y(_0888_));
 sky130_fd_sc_hd__clkinv_16 _1171_ (.A(net66),
    .Y(_0889_));
 sky130_fd_sc_hd__nand2_1 _1172_ (.A(net58),
    .B(net66),
    .Y(_0890_));
 sky130_fd_sc_hd__nand2_1 _1173_ (.A(net26),
    .B(net66),
    .Y(_0891_));
 sky130_fd_sc_hd__a21bo_1 _1174_ (.A1(sign),
    .A2(_0889_),
    .B1_N(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__mux2_1 _1175_ (.A0(_0874_),
    .A1(_0892_),
    .S(_0890_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _1176_ (.A0(\abs_multiplier[0] ),
    .A1(net34),
    .S(net66),
    .X(_0001_));
 sky130_fd_sc_hd__nand2_1 _1177_ (.A(net58),
    .B(net34),
    .Y(_0893_));
 sky130_fd_sc_hd__xnor2_1 _1178_ (.A(net45),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__mux2_1 _1179_ (.A0(\abs_multiplier[1] ),
    .A1(_0894_),
    .S(net66),
    .X(_0002_));
 sky130_fd_sc_hd__o21ai_1 _1180_ (.A1(net34),
    .A2(net45),
    .B1(net58),
    .Y(_0895_));
 sky130_fd_sc_hd__xnor2_1 _1181_ (.A(net56),
    .B(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__mux2_1 _1182_ (.A0(\abs_multiplier[2] ),
    .A1(_0896_),
    .S(net66),
    .X(_0003_));
 sky130_fd_sc_hd__o31a_1 _1183_ (.A1(net34),
    .A2(net45),
    .A3(net56),
    .B1(net58),
    .X(_0897_));
 sky130_fd_sc_hd__xor2_1 _1184_ (.A(net59),
    .B(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _1185_ (.A0(\abs_multiplier[3] ),
    .A1(_0898_),
    .S(net66),
    .X(_0004_));
 sky130_fd_sc_hd__or4_2 _1186_ (.A(net34),
    .B(net45),
    .C(net56),
    .D(net59),
    .X(_0899_));
 sky130_fd_sc_hd__a21oi_1 _1187_ (.A1(net58),
    .A2(_0899_),
    .B1(net60),
    .Y(_0900_));
 sky130_fd_sc_hd__a31o_1 _1188_ (.A1(net58),
    .A2(net60),
    .A3(_0899_),
    .B1(_0889_),
    .X(_0901_));
 sky130_fd_sc_hd__a2bb2o_1 _1189_ (.A1_N(_0900_),
    .A2_N(_0901_),
    .B1(\abs_multiplier[4] ),
    .B2(_0889_),
    .X(_0005_));
 sky130_fd_sc_hd__o21ai_1 _1190_ (.A1(net60),
    .A2(_0899_),
    .B1(net58),
    .Y(_0902_));
 sky130_fd_sc_hd__xnor2_1 _1191_ (.A(net61),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__mux2_1 _1192_ (.A0(\abs_multiplier[5] ),
    .A1(_0903_),
    .S(net66),
    .X(_0006_));
 sky130_fd_sc_hd__o31a_1 _1193_ (.A1(net60),
    .A2(net61),
    .A3(_0899_),
    .B1(net58),
    .X(_0904_));
 sky130_fd_sc_hd__xor2_1 _1194_ (.A(net62),
    .B(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__mux2_1 _1195_ (.A0(\abs_multiplier[6] ),
    .A1(_0905_),
    .S(net66),
    .X(_0007_));
 sky130_fd_sc_hd__or4_2 _1196_ (.A(net60),
    .B(net61),
    .C(net62),
    .D(_0899_),
    .X(_0906_));
 sky130_fd_sc_hd__a21oi_1 _1197_ (.A1(net58),
    .A2(_0906_),
    .B1(net63),
    .Y(_0907_));
 sky130_fd_sc_hd__a31o_1 _1198_ (.A1(net58),
    .A2(net63),
    .A3(_0906_),
    .B1(_0889_),
    .X(_0908_));
 sky130_fd_sc_hd__a2bb2o_1 _1199_ (.A1_N(_0907_),
    .A2_N(_0908_),
    .B1(\abs_multiplier[7] ),
    .B2(_0889_),
    .X(_0008_));
 sky130_fd_sc_hd__o21ai_1 _1200_ (.A1(net63),
    .A2(_0906_),
    .B1(net58),
    .Y(_0909_));
 sky130_fd_sc_hd__and2_1 _1201_ (.A(net64),
    .B(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__o21ai_1 _1202_ (.A1(net64),
    .A2(_0909_),
    .B1(net66),
    .Y(_0911_));
 sky130_fd_sc_hd__o22a_1 _1203_ (.A1(\abs_multiplier[8] ),
    .A2(net66),
    .B1(_0910_),
    .B2(_0911_),
    .X(_0009_));
 sky130_fd_sc_hd__or3_2 _1204_ (.A(net63),
    .B(net64),
    .C(_0906_),
    .X(_0912_));
 sky130_fd_sc_hd__a21oi_1 _1205_ (.A1(net58),
    .A2(_0912_),
    .B1(net65),
    .Y(_0913_));
 sky130_fd_sc_hd__a31o_1 _1206_ (.A1(net58),
    .A2(net65),
    .A3(_0912_),
    .B1(_0889_),
    .X(_0914_));
 sky130_fd_sc_hd__a2bb2o_1 _1207_ (.A1_N(_0913_),
    .A2_N(_0914_),
    .B1(\abs_multiplier[9] ),
    .B2(_0889_),
    .X(_0010_));
 sky130_fd_sc_hd__o21ai_1 _1208_ (.A1(net65),
    .A2(_0912_),
    .B1(net58),
    .Y(_0915_));
 sky130_fd_sc_hd__xnor2_1 _1209_ (.A(net35),
    .B(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__mux2_1 _1210_ (.A0(\abs_multiplier[10] ),
    .A1(_0916_),
    .S(net66),
    .X(_0011_));
 sky130_fd_sc_hd__o31a_1 _1211_ (.A1(net65),
    .A2(net35),
    .A3(_0912_),
    .B1(net58),
    .X(_0917_));
 sky130_fd_sc_hd__xor2_1 _1212_ (.A(net36),
    .B(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _1213_ (.A0(\abs_multiplier[11] ),
    .A1(_0918_),
    .S(net66),
    .X(_0012_));
 sky130_fd_sc_hd__or4_2 _1214_ (.A(net65),
    .B(net35),
    .C(net36),
    .D(_0912_),
    .X(_0919_));
 sky130_fd_sc_hd__a21oi_1 _1215_ (.A1(net58),
    .A2(_0919_),
    .B1(net37),
    .Y(_0920_));
 sky130_fd_sc_hd__a31o_1 _1216_ (.A1(net58),
    .A2(net37),
    .A3(_0919_),
    .B1(_0889_),
    .X(_0921_));
 sky130_fd_sc_hd__a2bb2o_1 _1217_ (.A1_N(_0920_),
    .A2_N(_0921_),
    .B1(\abs_multiplier[12] ),
    .B2(_0889_),
    .X(_0013_));
 sky130_fd_sc_hd__o21ai_1 _1218_ (.A1(net37),
    .A2(_0919_),
    .B1(net58),
    .Y(_0922_));
 sky130_fd_sc_hd__xnor2_1 _1219_ (.A(net38),
    .B(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__mux2_1 _1220_ (.A0(\abs_multiplier[13] ),
    .A1(_0923_),
    .S(net66),
    .X(_0014_));
 sky130_fd_sc_hd__or3_2 _1221_ (.A(net37),
    .B(net38),
    .C(_0919_),
    .X(_0924_));
 sky130_fd_sc_hd__a21oi_1 _1222_ (.A1(net58),
    .A2(_0924_),
    .B1(net39),
    .Y(_0925_));
 sky130_fd_sc_hd__a31o_1 _1223_ (.A1(net58),
    .A2(net39),
    .A3(_0924_),
    .B1(_0889_),
    .X(_0926_));
 sky130_fd_sc_hd__a2bb2o_1 _1224_ (.A1_N(_0925_),
    .A2_N(_0926_),
    .B1(\abs_multiplier[14] ),
    .B2(_0889_),
    .X(_0015_));
 sky130_fd_sc_hd__o21ai_1 _1225_ (.A1(net39),
    .A2(_0924_),
    .B1(net58),
    .Y(_0927_));
 sky130_fd_sc_hd__xnor2_1 _1226_ (.A(net40),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__mux2_1 _1227_ (.A0(\abs_multiplier[15] ),
    .A1(_0928_),
    .S(net66),
    .X(_0016_));
 sky130_fd_sc_hd__or3_1 _1228_ (.A(net39),
    .B(net40),
    .C(_0924_),
    .X(_0929_));
 sky130_fd_sc_hd__a21oi_1 _1229_ (.A1(net58),
    .A2(_0929_),
    .B1(_0886_),
    .Y(_0930_));
 sky130_fd_sc_hd__a31o_1 _1230_ (.A1(net58),
    .A2(_0886_),
    .A3(_0929_),
    .B1(_0889_),
    .X(_0931_));
 sky130_fd_sc_hd__o22a_1 _1231_ (.A1(\abs_multiplier[16] ),
    .A2(net66),
    .B1(_0930_),
    .B2(_0931_),
    .X(_0017_));
 sky130_fd_sc_hd__o21ai_1 _1232_ (.A1(net41),
    .A2(_0929_),
    .B1(net58),
    .Y(_0932_));
 sky130_fd_sc_hd__xnor2_1 _1233_ (.A(net42),
    .B(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__mux2_1 _1234_ (.A0(\abs_multiplier[17] ),
    .A1(_0933_),
    .S(net66),
    .X(_0018_));
 sky130_fd_sc_hd__or2_1 _1235_ (.A(net41),
    .B(net42),
    .X(_0934_));
 sky130_fd_sc_hd__or4_1 _1236_ (.A(net39),
    .B(net40),
    .C(_0924_),
    .D(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__a21oi_1 _1237_ (.A1(net58),
    .A2(_0935_),
    .B1(net43),
    .Y(_0936_));
 sky130_fd_sc_hd__a31o_1 _1238_ (.A1(net58),
    .A2(net43),
    .A3(_0935_),
    .B1(_0889_),
    .X(_0937_));
 sky130_fd_sc_hd__a2bb2o_1 _1239_ (.A1_N(_0936_),
    .A2_N(_0937_),
    .B1(\abs_multiplier[18] ),
    .B2(_0889_),
    .X(_0019_));
 sky130_fd_sc_hd__or2_1 _1240_ (.A(net43),
    .B(_0935_),
    .X(_0938_));
 sky130_fd_sc_hd__a21oi_1 _1241_ (.A1(net58),
    .A2(_0938_),
    .B1(net44),
    .Y(_0939_));
 sky130_fd_sc_hd__a31o_1 _1242_ (.A1(net58),
    .A2(net44),
    .A3(_0938_),
    .B1(_0889_),
    .X(_0940_));
 sky130_fd_sc_hd__a2bb2o_1 _1243_ (.A1_N(_0939_),
    .A2_N(_0940_),
    .B1(\abs_multiplier[19] ),
    .B2(_0889_),
    .X(_0020_));
 sky130_fd_sc_hd__or2_1 _1244_ (.A(net44),
    .B(_0938_),
    .X(_0941_));
 sky130_fd_sc_hd__a21oi_1 _1245_ (.A1(net58),
    .A2(_0941_),
    .B1(net46),
    .Y(_0942_));
 sky130_fd_sc_hd__a31o_1 _1246_ (.A1(net58),
    .A2(net46),
    .A3(_0941_),
    .B1(_0889_),
    .X(_0943_));
 sky130_fd_sc_hd__a2bb2o_1 _1247_ (.A1_N(_0942_),
    .A2_N(_0943_),
    .B1(\abs_multiplier[20] ),
    .B2(_0889_),
    .X(_0021_));
 sky130_fd_sc_hd__or3_1 _1248_ (.A(net44),
    .B(net46),
    .C(_0938_),
    .X(_0944_));
 sky130_fd_sc_hd__a21oi_1 _1249_ (.A1(net58),
    .A2(_0944_),
    .B1(net47),
    .Y(_0945_));
 sky130_fd_sc_hd__a31o_1 _1250_ (.A1(net58),
    .A2(net47),
    .A3(_0944_),
    .B1(_0889_),
    .X(_0946_));
 sky130_fd_sc_hd__a2bb2o_1 _1251_ (.A1_N(_0945_),
    .A2_N(_0946_),
    .B1(\abs_multiplier[21] ),
    .B2(_0889_),
    .X(_0022_));
 sky130_fd_sc_hd__o21ai_1 _1252_ (.A1(net47),
    .A2(_0944_),
    .B1(net58),
    .Y(_0947_));
 sky130_fd_sc_hd__xnor2_1 _1253_ (.A(net48),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__mux2_1 _1254_ (.A0(\abs_multiplier[22] ),
    .A1(_0948_),
    .S(net66),
    .X(_0023_));
 sky130_fd_sc_hd__or3_1 _1255_ (.A(net47),
    .B(net48),
    .C(_0944_),
    .X(_0949_));
 sky130_fd_sc_hd__a21oi_1 _1256_ (.A1(net58),
    .A2(_0949_),
    .B1(net49),
    .Y(_0950_));
 sky130_fd_sc_hd__a31o_1 _1257_ (.A1(net58),
    .A2(net49),
    .A3(_0949_),
    .B1(_0889_),
    .X(_0951_));
 sky130_fd_sc_hd__a2bb2o_1 _1258_ (.A1_N(_0950_),
    .A2_N(_0951_),
    .B1(\abs_multiplier[23] ),
    .B2(_0889_),
    .X(_0024_));
 sky130_fd_sc_hd__or2_2 _1259_ (.A(net49),
    .B(_0949_),
    .X(_0952_));
 sky130_fd_sc_hd__a21oi_1 _1260_ (.A1(net58),
    .A2(_0952_),
    .B1(_0887_),
    .Y(_0953_));
 sky130_fd_sc_hd__a31o_1 _1261_ (.A1(net58),
    .A2(_0887_),
    .A3(_0952_),
    .B1(_0889_),
    .X(_0954_));
 sky130_fd_sc_hd__o22a_1 _1262_ (.A1(\abs_multiplier[24] ),
    .A2(net66),
    .B1(_0953_),
    .B2(_0954_),
    .X(_0025_));
 sky130_fd_sc_hd__o21ai_1 _1263_ (.A1(net50),
    .A2(_0952_),
    .B1(net58),
    .Y(_0955_));
 sky130_fd_sc_hd__xnor2_1 _1264_ (.A(net51),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__mux2_1 _1265_ (.A0(\abs_multiplier[25] ),
    .A1(_0956_),
    .S(net66),
    .X(_0026_));
 sky130_fd_sc_hd__or2_1 _1266_ (.A(net50),
    .B(net51),
    .X(_0957_));
 sky130_fd_sc_hd__o21a_1 _1267_ (.A1(_0952_),
    .A2(_0957_),
    .B1(net58),
    .X(_0958_));
 sky130_fd_sc_hd__xor2_1 _1268_ (.A(net52),
    .B(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _1269_ (.A0(\abs_multiplier[26] ),
    .A1(_0959_),
    .S(net66),
    .X(_0027_));
 sky130_fd_sc_hd__o31a_1 _1270_ (.A1(net52),
    .A2(_0952_),
    .A3(_0957_),
    .B1(net58),
    .X(_0960_));
 sky130_fd_sc_hd__or2_1 _1271_ (.A(net53),
    .B(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__a21oi_1 _1272_ (.A1(net53),
    .A2(_0960_),
    .B1(_0889_),
    .Y(_0962_));
 sky130_fd_sc_hd__a22o_1 _1273_ (.A1(\abs_multiplier[27] ),
    .A2(_0889_),
    .B1(_0961_),
    .B2(_0962_),
    .X(_0028_));
 sky130_fd_sc_hd__or4_1 _1274_ (.A(net52),
    .B(net53),
    .C(_0952_),
    .D(_0957_),
    .X(_0963_));
 sky130_fd_sc_hd__nand2_1 _1275_ (.A(net58),
    .B(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__xnor2_1 _1276_ (.A(net54),
    .B(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__mux2_1 _1277_ (.A0(\abs_multiplier[28] ),
    .A1(_0965_),
    .S(net66),
    .X(_0029_));
 sky130_fd_sc_hd__or2_1 _1278_ (.A(net54),
    .B(_0963_),
    .X(_0966_));
 sky130_fd_sc_hd__a21oi_1 _1279_ (.A1(net58),
    .A2(_0966_),
    .B1(net55),
    .Y(_0967_));
 sky130_fd_sc_hd__a31o_1 _1280_ (.A1(net58),
    .A2(net55),
    .A3(_0966_),
    .B1(_0889_),
    .X(_0968_));
 sky130_fd_sc_hd__a2bb2o_1 _1281_ (.A1_N(_0967_),
    .A2_N(_0968_),
    .B1(\abs_multiplier[29] ),
    .B2(_0889_),
    .X(_0030_));
 sky130_fd_sc_hd__o21ai_1 _1282_ (.A1(net55),
    .A2(_0966_),
    .B1(net58),
    .Y(_0969_));
 sky130_fd_sc_hd__xnor2_1 _1283_ (.A(net57),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__mux2_1 _1284_ (.A0(\abs_multiplier[30] ),
    .A1(_0970_),
    .S(net66),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _1285_ (.A0(\abs_multiplicand[0] ),
    .A1(net2),
    .S(net66),
    .X(_0032_));
 sky130_fd_sc_hd__nand2_1 _1286_ (.A(net26),
    .B(net2),
    .Y(_0971_));
 sky130_fd_sc_hd__xnor2_1 _1287_ (.A(net13),
    .B(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__mux2_1 _1288_ (.A0(\abs_multiplicand[1] ),
    .A1(_0972_),
    .S(net66),
    .X(_0033_));
 sky130_fd_sc_hd__o21ai_1 _1289_ (.A1(net2),
    .A2(net13),
    .B1(net26),
    .Y(_0973_));
 sky130_fd_sc_hd__xnor2_1 _1290_ (.A(net24),
    .B(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__mux2_1 _1291_ (.A0(\abs_multiplicand[2] ),
    .A1(_0974_),
    .S(net66),
    .X(_0034_));
 sky130_fd_sc_hd__o31a_1 _1292_ (.A1(net2),
    .A2(net13),
    .A3(net24),
    .B1(net26),
    .X(_0975_));
 sky130_fd_sc_hd__xor2_1 _1293_ (.A(net27),
    .B(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__mux2_1 _1294_ (.A0(\abs_multiplicand[3] ),
    .A1(_0976_),
    .S(net66),
    .X(_0035_));
 sky130_fd_sc_hd__or4_2 _1295_ (.A(net2),
    .B(net13),
    .C(net24),
    .D(net27),
    .X(_0977_));
 sky130_fd_sc_hd__a21oi_1 _1296_ (.A1(net26),
    .A2(_0977_),
    .B1(net28),
    .Y(_0978_));
 sky130_fd_sc_hd__a31o_1 _1297_ (.A1(net26),
    .A2(net28),
    .A3(_0977_),
    .B1(_0889_),
    .X(_0979_));
 sky130_fd_sc_hd__a2bb2o_1 _1298_ (.A1_N(_0978_),
    .A2_N(_0979_),
    .B1(\abs_multiplicand[4] ),
    .B2(_0889_),
    .X(_0036_));
 sky130_fd_sc_hd__o21ai_1 _1299_ (.A1(net28),
    .A2(_0977_),
    .B1(net26),
    .Y(_0980_));
 sky130_fd_sc_hd__xnor2_1 _1300_ (.A(net29),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__mux2_1 _1301_ (.A0(\abs_multiplicand[5] ),
    .A1(_0981_),
    .S(net66),
    .X(_0037_));
 sky130_fd_sc_hd__o31a_1 _1302_ (.A1(net28),
    .A2(net29),
    .A3(_0977_),
    .B1(net26),
    .X(_0982_));
 sky130_fd_sc_hd__xor2_1 _1303_ (.A(net30),
    .B(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_1 _1304_ (.A0(\abs_multiplicand[6] ),
    .A1(_0983_),
    .S(net66),
    .X(_0038_));
 sky130_fd_sc_hd__or4_2 _1305_ (.A(net28),
    .B(net29),
    .C(net30),
    .D(_0977_),
    .X(_0984_));
 sky130_fd_sc_hd__a21oi_1 _1306_ (.A1(net26),
    .A2(_0984_),
    .B1(net31),
    .Y(_0985_));
 sky130_fd_sc_hd__a31o_1 _1307_ (.A1(net26),
    .A2(net31),
    .A3(_0984_),
    .B1(_0889_),
    .X(_0986_));
 sky130_fd_sc_hd__a2bb2o_1 _1308_ (.A1_N(_0985_),
    .A2_N(_0986_),
    .B1(\abs_multiplicand[7] ),
    .B2(_0889_),
    .X(_0039_));
 sky130_fd_sc_hd__o21ai_1 _1309_ (.A1(net31),
    .A2(_0984_),
    .B1(net26),
    .Y(_0987_));
 sky130_fd_sc_hd__o21ai_1 _1310_ (.A1(net32),
    .A2(_0987_),
    .B1(net66),
    .Y(_0988_));
 sky130_fd_sc_hd__a21o_1 _1311_ (.A1(net32),
    .A2(_0987_),
    .B1(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__o21a_1 _1312_ (.A1(\abs_multiplicand[8] ),
    .A2(net66),
    .B1(_0989_),
    .X(_0040_));
 sky130_fd_sc_hd__or3_2 _1313_ (.A(net31),
    .B(net32),
    .C(_0984_),
    .X(_0990_));
 sky130_fd_sc_hd__a21oi_1 _1314_ (.A1(net26),
    .A2(_0990_),
    .B1(net33),
    .Y(_0991_));
 sky130_fd_sc_hd__a31o_1 _1315_ (.A1(net26),
    .A2(net33),
    .A3(_0990_),
    .B1(_0889_),
    .X(_0992_));
 sky130_fd_sc_hd__a2bb2o_1 _1316_ (.A1_N(_0991_),
    .A2_N(_0992_),
    .B1(\abs_multiplicand[9] ),
    .B2(_0889_),
    .X(_0041_));
 sky130_fd_sc_hd__o21ai_1 _1317_ (.A1(net33),
    .A2(_0990_),
    .B1(net26),
    .Y(_0993_));
 sky130_fd_sc_hd__xnor2_1 _1318_ (.A(net3),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__mux2_1 _1319_ (.A0(\abs_multiplicand[10] ),
    .A1(_0994_),
    .S(net66),
    .X(_0042_));
 sky130_fd_sc_hd__o31a_1 _1320_ (.A1(net33),
    .A2(net3),
    .A3(_0990_),
    .B1(net26),
    .X(_0995_));
 sky130_fd_sc_hd__xor2_1 _1321_ (.A(net4),
    .B(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _1322_ (.A0(\abs_multiplicand[11] ),
    .A1(_0996_),
    .S(net66),
    .X(_0043_));
 sky130_fd_sc_hd__or4_1 _1323_ (.A(net33),
    .B(net3),
    .C(net4),
    .D(_0990_),
    .X(_0997_));
 sky130_fd_sc_hd__a21oi_1 _1324_ (.A1(net26),
    .A2(_0997_),
    .B1(net5),
    .Y(_0998_));
 sky130_fd_sc_hd__a31o_1 _1325_ (.A1(net26),
    .A2(net5),
    .A3(_0997_),
    .B1(_0889_),
    .X(_0999_));
 sky130_fd_sc_hd__a2bb2o_1 _1326_ (.A1_N(_0998_),
    .A2_N(_0999_),
    .B1(\abs_multiplicand[12] ),
    .B2(_0889_),
    .X(_0044_));
 sky130_fd_sc_hd__o21ai_1 _1327_ (.A1(net5),
    .A2(_0997_),
    .B1(net26),
    .Y(_1000_));
 sky130_fd_sc_hd__xnor2_1 _1328_ (.A(net6),
    .B(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__mux2_1 _1329_ (.A0(\abs_multiplicand[13] ),
    .A1(_1001_),
    .S(net66),
    .X(_0045_));
 sky130_fd_sc_hd__or3_1 _1330_ (.A(net5),
    .B(net6),
    .C(_0997_),
    .X(_1002_));
 sky130_fd_sc_hd__a21oi_1 _1331_ (.A1(net26),
    .A2(_1002_),
    .B1(net7),
    .Y(_1003_));
 sky130_fd_sc_hd__a31o_1 _1332_ (.A1(net26),
    .A2(net7),
    .A3(_1002_),
    .B1(_0889_),
    .X(_1004_));
 sky130_fd_sc_hd__a2bb2o_1 _1333_ (.A1_N(_1003_),
    .A2_N(_1004_),
    .B1(\abs_multiplicand[14] ),
    .B2(_0889_),
    .X(_0046_));
 sky130_fd_sc_hd__o21ai_1 _1334_ (.A1(net7),
    .A2(_1002_),
    .B1(net26),
    .Y(_1005_));
 sky130_fd_sc_hd__xnor2_1 _1335_ (.A(net8),
    .B(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__mux2_1 _1336_ (.A0(\abs_multiplicand[15] ),
    .A1(_1006_),
    .S(net66),
    .X(_0047_));
 sky130_fd_sc_hd__or3_2 _1337_ (.A(net7),
    .B(net8),
    .C(_1002_),
    .X(_1007_));
 sky130_fd_sc_hd__a21oi_1 _1338_ (.A1(net26),
    .A2(_1007_),
    .B1(_0884_),
    .Y(_1008_));
 sky130_fd_sc_hd__a31o_1 _1339_ (.A1(net26),
    .A2(_0884_),
    .A3(_1007_),
    .B1(_0889_),
    .X(_1009_));
 sky130_fd_sc_hd__o22a_1 _1340_ (.A1(\abs_multiplicand[16] ),
    .A2(net66),
    .B1(_1008_),
    .B2(_1009_),
    .X(_0048_));
 sky130_fd_sc_hd__o21ai_1 _1341_ (.A1(net9),
    .A2(_1007_),
    .B1(net26),
    .Y(_1010_));
 sky130_fd_sc_hd__xnor2_1 _1342_ (.A(net10),
    .B(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__mux2_1 _1343_ (.A0(\abs_multiplicand[17] ),
    .A1(_1011_),
    .S(net66),
    .X(_0049_));
 sky130_fd_sc_hd__o31a_1 _1344_ (.A1(net9),
    .A2(net10),
    .A3(_1007_),
    .B1(net26),
    .X(_1012_));
 sky130_fd_sc_hd__xor2_1 _1345_ (.A(net11),
    .B(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__mux2_1 _1346_ (.A0(\abs_multiplicand[18] ),
    .A1(_1013_),
    .S(net66),
    .X(_0050_));
 sky130_fd_sc_hd__or4_2 _1347_ (.A(net9),
    .B(net10),
    .C(net11),
    .D(_1007_),
    .X(_1014_));
 sky130_fd_sc_hd__a21oi_1 _1348_ (.A1(net26),
    .A2(_1014_),
    .B1(net12),
    .Y(_1015_));
 sky130_fd_sc_hd__a31o_1 _1349_ (.A1(net26),
    .A2(net12),
    .A3(_1014_),
    .B1(_0889_),
    .X(_1016_));
 sky130_fd_sc_hd__a2bb2o_1 _1350_ (.A1_N(_1015_),
    .A2_N(_1016_),
    .B1(\abs_multiplicand[19] ),
    .B2(_0889_),
    .X(_0051_));
 sky130_fd_sc_hd__o21ai_1 _1351_ (.A1(net12),
    .A2(_1014_),
    .B1(net26),
    .Y(_1017_));
 sky130_fd_sc_hd__xnor2_1 _1352_ (.A(net14),
    .B(_1017_),
    .Y(_1018_));
 sky130_fd_sc_hd__mux2_1 _1353_ (.A0(\abs_multiplicand[20] ),
    .A1(_1018_),
    .S(net66),
    .X(_0052_));
 sky130_fd_sc_hd__o31a_1 _1354_ (.A1(net12),
    .A2(net14),
    .A3(_1014_),
    .B1(net26),
    .X(_1019_));
 sky130_fd_sc_hd__xor2_1 _1355_ (.A(net15),
    .B(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(\abs_multiplicand[21] ),
    .A1(_1020_),
    .S(net66),
    .X(_0053_));
 sky130_fd_sc_hd__or4_1 _1357_ (.A(net12),
    .B(net14),
    .C(net15),
    .D(_1014_),
    .X(_1021_));
 sky130_fd_sc_hd__a21oi_1 _1358_ (.A1(net26),
    .A2(_1021_),
    .B1(net16),
    .Y(_1022_));
 sky130_fd_sc_hd__a31o_1 _1359_ (.A1(net26),
    .A2(net16),
    .A3(_1021_),
    .B1(_0889_),
    .X(_1023_));
 sky130_fd_sc_hd__a2bb2o_1 _1360_ (.A1_N(_1022_),
    .A2_N(_1023_),
    .B1(\abs_multiplicand[22] ),
    .B2(_0889_),
    .X(_0054_));
 sky130_fd_sc_hd__or2_1 _1361_ (.A(net16),
    .B(_1021_),
    .X(_1024_));
 sky130_fd_sc_hd__a21oi_1 _1362_ (.A1(net26),
    .A2(_1024_),
    .B1(net17),
    .Y(_1025_));
 sky130_fd_sc_hd__a31o_1 _1363_ (.A1(net26),
    .A2(net17),
    .A3(_1024_),
    .B1(_0889_),
    .X(_1026_));
 sky130_fd_sc_hd__a2bb2o_1 _1364_ (.A1_N(_1025_),
    .A2_N(_1026_),
    .B1(\abs_multiplicand[23] ),
    .B2(_0889_),
    .X(_0055_));
 sky130_fd_sc_hd__or2_1 _1365_ (.A(net17),
    .B(_1024_),
    .X(_1027_));
 sky130_fd_sc_hd__nand2_1 _1366_ (.A(net26),
    .B(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__o21ai_1 _1367_ (.A1(net18),
    .A2(_1028_),
    .B1(net66),
    .Y(_1029_));
 sky130_fd_sc_hd__a21o_1 _1368_ (.A1(net18),
    .A2(_1028_),
    .B1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__o21a_1 _1369_ (.A1(\abs_multiplicand[24] ),
    .A2(net66),
    .B1(_1030_),
    .X(_0056_));
 sky130_fd_sc_hd__o21ai_1 _1370_ (.A1(net18),
    .A2(_1027_),
    .B1(net26),
    .Y(_1031_));
 sky130_fd_sc_hd__xnor2_1 _1371_ (.A(net19),
    .B(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__mux2_1 _1372_ (.A0(\abs_multiplicand[25] ),
    .A1(_1032_),
    .S(net66),
    .X(_0057_));
 sky130_fd_sc_hd__o31a_1 _1373_ (.A1(net18),
    .A2(net19),
    .A3(_1027_),
    .B1(net26),
    .X(_1033_));
 sky130_fd_sc_hd__xor2_1 _1374_ (.A(net20),
    .B(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__mux2_1 _1375_ (.A0(\abs_multiplicand[26] ),
    .A1(_1034_),
    .S(net66),
    .X(_0058_));
 sky130_fd_sc_hd__or4_1 _1376_ (.A(net18),
    .B(net19),
    .C(net20),
    .D(_1027_),
    .X(_1035_));
 sky130_fd_sc_hd__a21oi_1 _1377_ (.A1(net26),
    .A2(_1035_),
    .B1(net21),
    .Y(_1036_));
 sky130_fd_sc_hd__a31o_1 _1378_ (.A1(net26),
    .A2(net21),
    .A3(_1035_),
    .B1(_0889_),
    .X(_1037_));
 sky130_fd_sc_hd__a2bb2o_1 _1379_ (.A1_N(_1036_),
    .A2_N(_1037_),
    .B1(\abs_multiplicand[27] ),
    .B2(_0889_),
    .X(_0059_));
 sky130_fd_sc_hd__or2_1 _1380_ (.A(net21),
    .B(_1035_),
    .X(_1038_));
 sky130_fd_sc_hd__a21oi_1 _1381_ (.A1(net26),
    .A2(_1038_),
    .B1(_0885_),
    .Y(_1039_));
 sky130_fd_sc_hd__a31o_1 _1382_ (.A1(net26),
    .A2(_0885_),
    .A3(_1038_),
    .B1(_0889_),
    .X(_1040_));
 sky130_fd_sc_hd__o22a_1 _1383_ (.A1(\abs_multiplicand[28] ),
    .A2(net66),
    .B1(_1039_),
    .B2(_1040_),
    .X(_0060_));
 sky130_fd_sc_hd__o21ai_1 _1384_ (.A1(net22),
    .A2(_1038_),
    .B1(net26),
    .Y(_1041_));
 sky130_fd_sc_hd__nor2_1 _1385_ (.A(net23),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__a21o_1 _1386_ (.A1(net23),
    .A2(_1041_),
    .B1(_0889_),
    .X(_1043_));
 sky130_fd_sc_hd__o22a_1 _1387_ (.A1(\abs_multiplicand[29] ),
    .A2(net66),
    .B1(_1042_),
    .B2(_1043_),
    .X(_0061_));
 sky130_fd_sc_hd__or3_1 _1388_ (.A(net22),
    .B(net23),
    .C(_1038_),
    .X(_1044_));
 sky130_fd_sc_hd__a21oi_1 _1389_ (.A1(net26),
    .A2(_1044_),
    .B1(net25),
    .Y(_1045_));
 sky130_fd_sc_hd__a31o_1 _1390_ (.A1(net26),
    .A2(net25),
    .A3(_1044_),
    .B1(_0889_),
    .X(_1046_));
 sky130_fd_sc_hd__a2bb2o_1 _1391_ (.A1_N(_1045_),
    .A2_N(_1046_),
    .B1(\abs_multiplicand[30] ),
    .B2(_0889_),
    .X(_0062_));
 sky130_fd_sc_hd__or2_2 _1392_ (.A(net135),
    .B(\count[4] ),
    .X(_1047_));
 sky130_fd_sc_hd__or4_4 _1393_ (.A(\count[3] ),
    .B(\count[2] ),
    .C(\count[1] ),
    .D(\count[0] ),
    .X(_1048_));
 sky130_fd_sc_hd__nor2_8 _1394_ (.A(_1047_),
    .B(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__or2_2 _1395_ (.A(_1047_),
    .B(_1048_),
    .X(_1050_));
 sky130_fd_sc_hd__mux2_1 _1396_ (.A0(\M[0] ),
    .A1(\abs_multiplicand[0] ),
    .S(_1049_),
    .X(_1051_));
 sky130_fd_sc_hd__and2_1 _1397_ (.A(_0889_),
    .B(_1051_),
    .X(_0063_));
 sky130_fd_sc_hd__or4b_1 _1398_ (.A(net135),
    .B(_1048_),
    .C(\count[4] ),
    .D_N(\abs_multiplicand[1] ),
    .X(_1052_));
 sky130_fd_sc_hd__or3_1 _1399_ (.A(\abs_multiplicand[1] ),
    .B(_1047_),
    .C(_1048_),
    .X(_1053_));
 sky130_fd_sc_hd__o21ai_1 _1400_ (.A1(_0883_),
    .A2(_1049_),
    .B1(_1052_),
    .Y(_1054_));
 sky130_fd_sc_hd__and2_1 _1401_ (.A(_0889_),
    .B(_1054_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1402_ (.A0(\M[2] ),
    .A1(\abs_multiplicand[2] ),
    .S(_1049_),
    .X(_1055_));
 sky130_fd_sc_hd__and2_1 _1403_ (.A(_0889_),
    .B(_1055_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1404_ (.A0(\M[3] ),
    .A1(\abs_multiplicand[3] ),
    .S(_1049_),
    .X(_1056_));
 sky130_fd_sc_hd__and2_1 _1405_ (.A(_0889_),
    .B(_1056_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1406_ (.A0(\M[4] ),
    .A1(\abs_multiplicand[4] ),
    .S(_1049_),
    .X(_1057_));
 sky130_fd_sc_hd__and2_1 _1407_ (.A(_0889_),
    .B(_1057_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1408_ (.A0(\M[5] ),
    .A1(\abs_multiplicand[5] ),
    .S(_1049_),
    .X(_1058_));
 sky130_fd_sc_hd__and2_1 _1409_ (.A(_0889_),
    .B(_1058_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1410_ (.A0(\M[6] ),
    .A1(\abs_multiplicand[6] ),
    .S(_1049_),
    .X(_1059_));
 sky130_fd_sc_hd__and2_1 _1411_ (.A(_0889_),
    .B(_1059_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_2 _1412_ (.A0(\M[7] ),
    .A1(\abs_multiplicand[7] ),
    .S(_1049_),
    .X(_1060_));
 sky130_fd_sc_hd__and2_1 _1413_ (.A(_0889_),
    .B(_1060_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1414_ (.A0(\M[8] ),
    .A1(\abs_multiplicand[8] ),
    .S(_1049_),
    .X(_1061_));
 sky130_fd_sc_hd__and2_1 _1415_ (.A(_0889_),
    .B(_1061_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1416_ (.A0(\M[9] ),
    .A1(\abs_multiplicand[9] ),
    .S(_1049_),
    .X(_1062_));
 sky130_fd_sc_hd__and2_1 _1417_ (.A(_0889_),
    .B(_1062_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1418_ (.A0(\M[10] ),
    .A1(\abs_multiplicand[10] ),
    .S(_1049_),
    .X(_1063_));
 sky130_fd_sc_hd__and2_1 _1419_ (.A(_0889_),
    .B(_1063_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1420_ (.A0(\M[11] ),
    .A1(\abs_multiplicand[11] ),
    .S(_1049_),
    .X(_1064_));
 sky130_fd_sc_hd__and2_1 _1421_ (.A(_0889_),
    .B(_1064_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1422_ (.A0(\M[12] ),
    .A1(\abs_multiplicand[12] ),
    .S(_1049_),
    .X(_1065_));
 sky130_fd_sc_hd__and2_1 _1423_ (.A(_0889_),
    .B(_1065_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_2 _1424_ (.A0(\M[13] ),
    .A1(\abs_multiplicand[13] ),
    .S(_1049_),
    .X(_1066_));
 sky130_fd_sc_hd__and2_1 _1425_ (.A(_0889_),
    .B(_1066_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1426_ (.A0(\M[14] ),
    .A1(\abs_multiplicand[14] ),
    .S(_1049_),
    .X(_1067_));
 sky130_fd_sc_hd__and2_1 _1427_ (.A(_0889_),
    .B(_1067_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1428_ (.A0(\M[15] ),
    .A1(\abs_multiplicand[15] ),
    .S(_1049_),
    .X(_1068_));
 sky130_fd_sc_hd__and2_1 _1429_ (.A(_0889_),
    .B(_1068_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _1430_ (.A0(\M[16] ),
    .A1(\abs_multiplicand[16] ),
    .S(net133),
    .X(_1069_));
 sky130_fd_sc_hd__and2_1 _1431_ (.A(_0889_),
    .B(_1069_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _1432_ (.A0(\M[17] ),
    .A1(\abs_multiplicand[17] ),
    .S(net133),
    .X(_1070_));
 sky130_fd_sc_hd__and2_1 _1433_ (.A(_0889_),
    .B(_1070_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1434_ (.A0(\M[18] ),
    .A1(\abs_multiplicand[18] ),
    .S(net133),
    .X(_1071_));
 sky130_fd_sc_hd__and2_1 _1435_ (.A(_0889_),
    .B(_1071_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _1436_ (.A0(\M[19] ),
    .A1(\abs_multiplicand[19] ),
    .S(net133),
    .X(_1072_));
 sky130_fd_sc_hd__and2_1 _1437_ (.A(_0889_),
    .B(_1072_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _1438_ (.A0(\M[20] ),
    .A1(\abs_multiplicand[20] ),
    .S(net133),
    .X(_1073_));
 sky130_fd_sc_hd__and2_1 _1439_ (.A(_0889_),
    .B(_1073_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(\M[21] ),
    .A1(\abs_multiplicand[21] ),
    .S(net133),
    .X(_1074_));
 sky130_fd_sc_hd__and2_1 _1441_ (.A(_0889_),
    .B(_1074_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _1442_ (.A0(\M[22] ),
    .A1(\abs_multiplicand[22] ),
    .S(net133),
    .X(_1075_));
 sky130_fd_sc_hd__and2_1 _1443_ (.A(_0889_),
    .B(_1075_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(\M[23] ),
    .A1(\abs_multiplicand[23] ),
    .S(net133),
    .X(_1076_));
 sky130_fd_sc_hd__and2_1 _1445_ (.A(_0889_),
    .B(_1076_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _1446_ (.A0(\M[24] ),
    .A1(\abs_multiplicand[24] ),
    .S(net133),
    .X(_1077_));
 sky130_fd_sc_hd__and2_1 _1447_ (.A(_0889_),
    .B(_1077_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _1448_ (.A0(\M[25] ),
    .A1(\abs_multiplicand[25] ),
    .S(net133),
    .X(_1078_));
 sky130_fd_sc_hd__and2_1 _1449_ (.A(_0889_),
    .B(_1078_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _1450_ (.A0(\M[26] ),
    .A1(\abs_multiplicand[26] ),
    .S(net133),
    .X(_1079_));
 sky130_fd_sc_hd__and2_1 _1451_ (.A(_0889_),
    .B(_1079_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1452_ (.A0(\M[27] ),
    .A1(\abs_multiplicand[27] ),
    .S(net133),
    .X(_1080_));
 sky130_fd_sc_hd__and2_1 _1453_ (.A(_0889_),
    .B(_1080_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _1454_ (.A0(\M[28] ),
    .A1(\abs_multiplicand[28] ),
    .S(net133),
    .X(_1081_));
 sky130_fd_sc_hd__and2_1 _1455_ (.A(_0889_),
    .B(_1081_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _1456_ (.A0(\M[29] ),
    .A1(\abs_multiplicand[29] ),
    .S(net133),
    .X(_1082_));
 sky130_fd_sc_hd__and2_1 _1457_ (.A(_0889_),
    .B(_1082_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _1458_ (.A0(\M[30] ),
    .A1(\abs_multiplicand[30] ),
    .S(net133),
    .X(_1083_));
 sky130_fd_sc_hd__and2_1 _1459_ (.A(_0889_),
    .B(_1083_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1460_ (.A0(\M[31] ),
    .A1(\abs_multiplicand[31] ),
    .S(net133),
    .X(_1084_));
 sky130_fd_sc_hd__and2_1 _1461_ (.A(_0889_),
    .B(_1084_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _1462_ (.A0(\Q[1] ),
    .A1(\abs_multiplier[1] ),
    .S(_1049_),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_1 _1463_ (.A0(\Q[0] ),
    .A1(_1085_),
    .S(_0873_),
    .X(_1086_));
 sky130_fd_sc_hd__and2_1 _1464_ (.A(_0889_),
    .B(_1086_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _1465_ (.A0(\Q[2] ),
    .A1(\abs_multiplier[2] ),
    .S(_1049_),
    .X(_1087_));
 sky130_fd_sc_hd__or2_1 _1466_ (.A(_0873_),
    .B(\Q[1] ),
    .X(_1088_));
 sky130_fd_sc_hd__o211a_1 _1467_ (.A1(net135),
    .A2(_1087_),
    .B1(_1088_),
    .C1(_0889_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _1468_ (.A0(\Q[3] ),
    .A1(\abs_multiplier[3] ),
    .S(_1049_),
    .X(_1089_));
 sky130_fd_sc_hd__or2_1 _1469_ (.A(_0873_),
    .B(\Q[2] ),
    .X(_1090_));
 sky130_fd_sc_hd__o211a_1 _1470_ (.A1(net135),
    .A2(_1089_),
    .B1(_1090_),
    .C1(_0889_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _1471_ (.A0(\Q[4] ),
    .A1(\abs_multiplier[4] ),
    .S(_1049_),
    .X(_1091_));
 sky130_fd_sc_hd__or2_1 _1472_ (.A(_0873_),
    .B(\Q[3] ),
    .X(_1092_));
 sky130_fd_sc_hd__o211a_1 _1473_ (.A1(net135),
    .A2(_1091_),
    .B1(_1092_),
    .C1(_0889_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _1474_ (.A0(\Q[5] ),
    .A1(\abs_multiplier[5] ),
    .S(_1049_),
    .X(_1093_));
 sky130_fd_sc_hd__nand2_1 _1475_ (.A(net135),
    .B(_0882_),
    .Y(_1094_));
 sky130_fd_sc_hd__o211a_1 _1476_ (.A1(net135),
    .A2(_1093_),
    .B1(_1094_),
    .C1(_0889_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(\Q[6] ),
    .A1(\abs_multiplier[6] ),
    .S(_1049_),
    .X(_1095_));
 sky130_fd_sc_hd__or2_1 _1478_ (.A(_0873_),
    .B(\Q[5] ),
    .X(_1096_));
 sky130_fd_sc_hd__o211a_1 _1479_ (.A1(net135),
    .A2(_1095_),
    .B1(_1096_),
    .C1(_0889_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _1480_ (.A0(\Q[7] ),
    .A1(\abs_multiplier[7] ),
    .S(_1049_),
    .X(_1097_));
 sky130_fd_sc_hd__or2_1 _1481_ (.A(_0873_),
    .B(\Q[6] ),
    .X(_1098_));
 sky130_fd_sc_hd__o211a_1 _1482_ (.A1(net135),
    .A2(_1097_),
    .B1(_1098_),
    .C1(_0889_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1483_ (.A0(\Q[8] ),
    .A1(\abs_multiplier[8] ),
    .S(_1049_),
    .X(_1099_));
 sky130_fd_sc_hd__or2_1 _1484_ (.A(_0873_),
    .B(\Q[7] ),
    .X(_1100_));
 sky130_fd_sc_hd__o211a_1 _1485_ (.A1(net135),
    .A2(_1099_),
    .B1(_1100_),
    .C1(_0889_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(\Q[9] ),
    .A1(\abs_multiplier[9] ),
    .S(_1049_),
    .X(_1101_));
 sky130_fd_sc_hd__or2_1 _1487_ (.A(_0873_),
    .B(\Q[8] ),
    .X(_1102_));
 sky130_fd_sc_hd__o211a_1 _1488_ (.A1(net135),
    .A2(_1101_),
    .B1(_1102_),
    .C1(_0889_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1489_ (.A0(\Q[10] ),
    .A1(\abs_multiplier[10] ),
    .S(_1049_),
    .X(_1103_));
 sky130_fd_sc_hd__or2_1 _1490_ (.A(_0873_),
    .B(\Q[9] ),
    .X(_1104_));
 sky130_fd_sc_hd__o211a_1 _1491_ (.A1(net135),
    .A2(_1103_),
    .B1(_1104_),
    .C1(_0889_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1492_ (.A0(\Q[11] ),
    .A1(\abs_multiplier[11] ),
    .S(net133),
    .X(_1105_));
 sky130_fd_sc_hd__nand2_1 _1493_ (.A(net135),
    .B(_0881_),
    .Y(_1106_));
 sky130_fd_sc_hd__o211a_1 _1494_ (.A1(net135),
    .A2(_1105_),
    .B1(_1106_),
    .C1(_0889_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(\Q[12] ),
    .A1(\abs_multiplier[12] ),
    .S(net133),
    .X(_1107_));
 sky130_fd_sc_hd__or2_1 _1496_ (.A(_0873_),
    .B(\Q[11] ),
    .X(_1108_));
 sky130_fd_sc_hd__o211a_1 _1497_ (.A1(net135),
    .A2(_1107_),
    .B1(_1108_),
    .C1(_0889_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1498_ (.A0(\Q[13] ),
    .A1(\abs_multiplier[13] ),
    .S(net133),
    .X(_1109_));
 sky130_fd_sc_hd__or2_1 _1499_ (.A(_0873_),
    .B(\Q[12] ),
    .X(_1110_));
 sky130_fd_sc_hd__o211a_1 _1500_ (.A1(net135),
    .A2(_1109_),
    .B1(_1110_),
    .C1(_0889_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1501_ (.A0(\Q[14] ),
    .A1(\abs_multiplier[14] ),
    .S(net133),
    .X(_1111_));
 sky130_fd_sc_hd__nand2_1 _1502_ (.A(net134),
    .B(_0880_),
    .Y(_1112_));
 sky130_fd_sc_hd__o211a_1 _1503_ (.A1(net134),
    .A2(_1111_),
    .B1(_1112_),
    .C1(_0889_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1504_ (.A0(\Q[15] ),
    .A1(\abs_multiplier[15] ),
    .S(net133),
    .X(_1113_));
 sky130_fd_sc_hd__or2_1 _1505_ (.A(_0873_),
    .B(\Q[14] ),
    .X(_1114_));
 sky130_fd_sc_hd__o211a_1 _1506_ (.A1(net134),
    .A2(_1113_),
    .B1(_1114_),
    .C1(_0889_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1507_ (.A0(\Q[16] ),
    .A1(\abs_multiplier[16] ),
    .S(net133),
    .X(_1115_));
 sky130_fd_sc_hd__or2_1 _1508_ (.A(_0873_),
    .B(\Q[15] ),
    .X(_1116_));
 sky130_fd_sc_hd__o211a_1 _1509_ (.A1(net134),
    .A2(_1115_),
    .B1(_1116_),
    .C1(_0889_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _1510_ (.A0(\Q[17] ),
    .A1(\abs_multiplier[17] ),
    .S(net133),
    .X(_1117_));
 sky130_fd_sc_hd__or2_1 _1511_ (.A(_0873_),
    .B(\Q[16] ),
    .X(_1118_));
 sky130_fd_sc_hd__o211a_1 _1512_ (.A1(net134),
    .A2(_1117_),
    .B1(_1118_),
    .C1(_0889_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _1513_ (.A0(\Q[18] ),
    .A1(\abs_multiplier[18] ),
    .S(net133),
    .X(_1119_));
 sky130_fd_sc_hd__or2_1 _1514_ (.A(_0873_),
    .B(\Q[17] ),
    .X(_1120_));
 sky130_fd_sc_hd__o211a_1 _1515_ (.A1(net134),
    .A2(_1119_),
    .B1(_1120_),
    .C1(_0889_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1516_ (.A0(\Q[19] ),
    .A1(\abs_multiplier[19] ),
    .S(net133),
    .X(_1121_));
 sky130_fd_sc_hd__or2_1 _1517_ (.A(_0873_),
    .B(\Q[18] ),
    .X(_1122_));
 sky130_fd_sc_hd__o211a_1 _1518_ (.A1(net134),
    .A2(_1121_),
    .B1(_1122_),
    .C1(_0889_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1519_ (.A0(\Q[20] ),
    .A1(\abs_multiplier[20] ),
    .S(net133),
    .X(_1123_));
 sky130_fd_sc_hd__or2_1 _1520_ (.A(_0873_),
    .B(\Q[19] ),
    .X(_1124_));
 sky130_fd_sc_hd__o211a_1 _1521_ (.A1(net134),
    .A2(_1123_),
    .B1(_1124_),
    .C1(_0889_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1522_ (.A0(\Q[21] ),
    .A1(\abs_multiplier[21] ),
    .S(net133),
    .X(_1125_));
 sky130_fd_sc_hd__or2_1 _1523_ (.A(_0873_),
    .B(\Q[20] ),
    .X(_1126_));
 sky130_fd_sc_hd__o211a_1 _1524_ (.A1(net134),
    .A2(_1125_),
    .B1(_1126_),
    .C1(_0889_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _1525_ (.A0(\Q[22] ),
    .A1(\abs_multiplier[22] ),
    .S(net133),
    .X(_1127_));
 sky130_fd_sc_hd__or2_1 _1526_ (.A(_0873_),
    .B(\Q[21] ),
    .X(_1128_));
 sky130_fd_sc_hd__o211a_1 _1527_ (.A1(net134),
    .A2(_1127_),
    .B1(_1128_),
    .C1(_0889_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _1528_ (.A0(\Q[23] ),
    .A1(\abs_multiplier[23] ),
    .S(net133),
    .X(_1129_));
 sky130_fd_sc_hd__nand2_1 _1529_ (.A(net134),
    .B(_0879_),
    .Y(_1130_));
 sky130_fd_sc_hd__o211a_1 _1530_ (.A1(net134),
    .A2(_1129_),
    .B1(_1130_),
    .C1(_0889_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1531_ (.A0(\Q[24] ),
    .A1(\abs_multiplier[24] ),
    .S(net133),
    .X(_1131_));
 sky130_fd_sc_hd__or2_1 _1532_ (.A(_0873_),
    .B(\Q[23] ),
    .X(_1132_));
 sky130_fd_sc_hd__o211a_1 _1533_ (.A1(net134),
    .A2(_1131_),
    .B1(_1132_),
    .C1(_0889_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _1534_ (.A0(\Q[25] ),
    .A1(\abs_multiplier[25] ),
    .S(net133),
    .X(_1133_));
 sky130_fd_sc_hd__nand2_1 _1535_ (.A(net134),
    .B(_0878_),
    .Y(_1134_));
 sky130_fd_sc_hd__o211a_1 _1536_ (.A1(net134),
    .A2(_1133_),
    .B1(_1134_),
    .C1(_0889_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _1537_ (.A0(\Q[26] ),
    .A1(\abs_multiplier[26] ),
    .S(net133),
    .X(_1135_));
 sky130_fd_sc_hd__or2_1 _1538_ (.A(_0873_),
    .B(\Q[25] ),
    .X(_1136_));
 sky130_fd_sc_hd__o211a_1 _1539_ (.A1(net134),
    .A2(_1135_),
    .B1(_1136_),
    .C1(_0889_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _1540_ (.A0(\Q[27] ),
    .A1(\abs_multiplier[27] ),
    .S(net133),
    .X(_1137_));
 sky130_fd_sc_hd__or2_1 _1541_ (.A(_0873_),
    .B(\Q[26] ),
    .X(_1138_));
 sky130_fd_sc_hd__o211a_1 _1542_ (.A1(net134),
    .A2(_1137_),
    .B1(_1138_),
    .C1(_0889_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _1543_ (.A0(\Q[28] ),
    .A1(\abs_multiplier[28] ),
    .S(net133),
    .X(_1139_));
 sky130_fd_sc_hd__or2_1 _1544_ (.A(_0873_),
    .B(\Q[27] ),
    .X(_1140_));
 sky130_fd_sc_hd__o211a_1 _1545_ (.A1(net134),
    .A2(_1139_),
    .B1(_1140_),
    .C1(_0889_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1546_ (.A0(\Q[29] ),
    .A1(\abs_multiplier[29] ),
    .S(net133),
    .X(_1141_));
 sky130_fd_sc_hd__nand2_1 _1547_ (.A(net135),
    .B(_0877_),
    .Y(_1142_));
 sky130_fd_sc_hd__o211a_1 _1548_ (.A1(net135),
    .A2(_1141_),
    .B1(_1142_),
    .C1(_0889_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1549_ (.A0(\Q[30] ),
    .A1(\abs_multiplier[30] ),
    .S(net133),
    .X(_1143_));
 sky130_fd_sc_hd__or2_1 _1550_ (.A(_0873_),
    .B(\Q[29] ),
    .X(_1144_));
 sky130_fd_sc_hd__o211a_1 _1551_ (.A1(net135),
    .A2(_1143_),
    .B1(_1144_),
    .C1(_0889_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(\Q[31] ),
    .A1(\abs_multiplier[31] ),
    .S(net133),
    .X(_1145_));
 sky130_fd_sc_hd__or2_1 _1553_ (.A(net135),
    .B(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__o211a_1 _1554_ (.A1(_0873_),
    .A2(\Q[30] ),
    .B1(_0889_),
    .C1(_1146_),
    .X(_0125_));
 sky130_fd_sc_hd__or2_1 _1555_ (.A(\Q[0] ),
    .B(_1049_),
    .X(_1147_));
 sky130_fd_sc_hd__o21a_4 _1556_ (.A1(\abs_multiplier[0] ),
    .A2(_1050_),
    .B1(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__o21ai_4 _1557_ (.A1(\abs_multiplier[0] ),
    .A2(_1050_),
    .B1(_1147_),
    .Y(_1149_));
 sky130_fd_sc_hd__nand2_1 _1558_ (.A(_1051_),
    .B(_1148_),
    .Y(_1150_));
 sky130_fd_sc_hd__xnor2_1 _1559_ (.A(\A[0] ),
    .B(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__or2_1 _1560_ (.A(_0873_),
    .B(\Q[31] ),
    .X(_0263_));
 sky130_fd_sc_hd__o211a_1 _1561_ (.A1(net135),
    .A2(_1151_),
    .B1(_0263_),
    .C1(_0889_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1562_ (.A0(net68),
    .A1(\Q[0] ),
    .S(net135),
    .X(_0264_));
 sky130_fd_sc_hd__and2_1 _1563_ (.A(_0889_),
    .B(_0264_),
    .X(_0127_));
 sky130_fd_sc_hd__and3_1 _1564_ (.A(\Q[0] ),
    .B(\Q[1] ),
    .C(sign),
    .X(_0265_));
 sky130_fd_sc_hd__a21oi_1 _1565_ (.A1(\Q[0] ),
    .A2(sign),
    .B1(\Q[1] ),
    .Y(_0266_));
 sky130_fd_sc_hd__o21ai_1 _1566_ (.A1(_0265_),
    .A2(_0266_),
    .B1(net135),
    .Y(_0267_));
 sky130_fd_sc_hd__o211a_1 _1567_ (.A1(net135),
    .A2(net79),
    .B1(_0889_),
    .C1(_0267_),
    .X(_0128_));
 sky130_fd_sc_hd__o21ai_1 _1568_ (.A1(\Q[0] ),
    .A2(\Q[1] ),
    .B1(sign),
    .Y(_0268_));
 sky130_fd_sc_hd__nor2_1 _1569_ (.A(\Q[2] ),
    .B(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__and2_1 _1570_ (.A(\Q[2] ),
    .B(_0268_),
    .X(_0270_));
 sky130_fd_sc_hd__or2_1 _1571_ (.A(net135),
    .B(net90),
    .X(_0271_));
 sky130_fd_sc_hd__o311a_1 _1572_ (.A1(_0873_),
    .A2(_0269_),
    .A3(_0270_),
    .B1(_0271_),
    .C1(_0889_),
    .X(_0129_));
 sky130_fd_sc_hd__o31a_1 _1573_ (.A1(\Q[0] ),
    .A2(\Q[2] ),
    .A3(\Q[1] ),
    .B1(sign),
    .X(_0272_));
 sky130_fd_sc_hd__xor2_1 _1574_ (.A(\Q[3] ),
    .B(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__or2_1 _1575_ (.A(net135),
    .B(net101),
    .X(_0274_));
 sky130_fd_sc_hd__o211a_1 _1576_ (.A1(_0873_),
    .A2(_0273_),
    .B1(_0274_),
    .C1(_0889_),
    .X(_0130_));
 sky130_fd_sc_hd__or4_2 _1577_ (.A(\Q[0] ),
    .B(\Q[3] ),
    .C(\Q[2] ),
    .D(\Q[1] ),
    .X(_0275_));
 sky130_fd_sc_hd__a21oi_1 _1578_ (.A1(sign),
    .A2(_0275_),
    .B1(_0882_),
    .Y(_0276_));
 sky130_fd_sc_hd__a31o_1 _1579_ (.A1(_0882_),
    .A2(sign),
    .A3(_0275_),
    .B1(_0873_),
    .X(_0277_));
 sky130_fd_sc_hd__o221a_1 _1580_ (.A1(net135),
    .A2(net112),
    .B1(_0276_),
    .B2(_0277_),
    .C1(_0889_),
    .X(_0131_));
 sky130_fd_sc_hd__o21ai_1 _1581_ (.A1(\Q[4] ),
    .A2(_0275_),
    .B1(sign),
    .Y(_0278_));
 sky130_fd_sc_hd__xnor2_1 _1582_ (.A(\Q[5] ),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__or2_1 _1583_ (.A(net135),
    .B(net123),
    .X(_0280_));
 sky130_fd_sc_hd__o211a_1 _1584_ (.A1(_0873_),
    .A2(_0279_),
    .B1(_0280_),
    .C1(_0889_),
    .X(_0132_));
 sky130_fd_sc_hd__o31a_1 _1585_ (.A1(\Q[5] ),
    .A2(\Q[4] ),
    .A3(_0275_),
    .B1(sign),
    .X(_0281_));
 sky130_fd_sc_hd__xor2_1 _1586_ (.A(\Q[6] ),
    .B(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__or2_1 _1587_ (.A(net135),
    .B(net128),
    .X(_0283_));
 sky130_fd_sc_hd__o211a_1 _1588_ (.A1(_0873_),
    .A2(_0282_),
    .B1(_0283_),
    .C1(_0889_),
    .X(_0133_));
 sky130_fd_sc_hd__or4_2 _1589_ (.A(\Q[6] ),
    .B(\Q[5] ),
    .C(\Q[4] ),
    .D(_0275_),
    .X(_0284_));
 sky130_fd_sc_hd__and3_1 _1590_ (.A(\Q[7] ),
    .B(sign),
    .C(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__a21oi_1 _1591_ (.A1(sign),
    .A2(_0284_),
    .B1(\Q[7] ),
    .Y(_0286_));
 sky130_fd_sc_hd__o21ai_1 _1592_ (.A1(_0285_),
    .A2(_0286_),
    .B1(net135),
    .Y(_0287_));
 sky130_fd_sc_hd__o211a_1 _1593_ (.A1(net135),
    .A2(net129),
    .B1(_0889_),
    .C1(_0287_),
    .X(_0134_));
 sky130_fd_sc_hd__o21ai_1 _1594_ (.A1(\Q[7] ),
    .A2(_0284_),
    .B1(sign),
    .Y(_0288_));
 sky130_fd_sc_hd__xnor2_1 _1595_ (.A(\Q[8] ),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__or2_1 _1596_ (.A(net135),
    .B(net130),
    .X(_0290_));
 sky130_fd_sc_hd__o211a_1 _1597_ (.A1(_0873_),
    .A2(_0289_),
    .B1(_0290_),
    .C1(_0889_),
    .X(_0135_));
 sky130_fd_sc_hd__o31a_1 _1598_ (.A1(\Q[8] ),
    .A2(\Q[7] ),
    .A3(_0284_),
    .B1(sign),
    .X(_0291_));
 sky130_fd_sc_hd__xor2_1 _1599_ (.A(\Q[9] ),
    .B(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _1600_ (.A(net135),
    .B(net131),
    .X(_0293_));
 sky130_fd_sc_hd__o211a_1 _1601_ (.A1(_0873_),
    .A2(_0292_),
    .B1(_0293_),
    .C1(_0889_),
    .X(_0136_));
 sky130_fd_sc_hd__or4_2 _1602_ (.A(\Q[9] ),
    .B(\Q[8] ),
    .C(\Q[7] ),
    .D(_0284_),
    .X(_0294_));
 sky130_fd_sc_hd__and3_1 _1603_ (.A(_0881_),
    .B(sign),
    .C(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__a21oi_1 _1604_ (.A1(sign),
    .A2(_0294_),
    .B1(_0881_),
    .Y(_0296_));
 sky130_fd_sc_hd__or2_1 _1605_ (.A(net135),
    .B(net69),
    .X(_0297_));
 sky130_fd_sc_hd__o311a_1 _1606_ (.A1(_0873_),
    .A2(_0295_),
    .A3(_0296_),
    .B1(_0297_),
    .C1(_0889_),
    .X(_0137_));
 sky130_fd_sc_hd__o21ai_1 _1607_ (.A1(\Q[10] ),
    .A2(_0294_),
    .B1(sign),
    .Y(_0298_));
 sky130_fd_sc_hd__xnor2_1 _1608_ (.A(\Q[11] ),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__or2_1 _1609_ (.A(net135),
    .B(net70),
    .X(_0300_));
 sky130_fd_sc_hd__o211a_1 _1610_ (.A1(_0873_),
    .A2(_0299_),
    .B1(_0300_),
    .C1(_0889_),
    .X(_0138_));
 sky130_fd_sc_hd__o31a_1 _1611_ (.A1(\Q[11] ),
    .A2(\Q[10] ),
    .A3(_0294_),
    .B1(sign),
    .X(_0301_));
 sky130_fd_sc_hd__xor2_1 _1612_ (.A(\Q[12] ),
    .B(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__or2_1 _1613_ (.A(net135),
    .B(net71),
    .X(_0303_));
 sky130_fd_sc_hd__o211a_1 _1614_ (.A1(_0873_),
    .A2(_0302_),
    .B1(_0303_),
    .C1(_0889_),
    .X(_0139_));
 sky130_fd_sc_hd__or4_2 _1615_ (.A(\Q[12] ),
    .B(\Q[11] ),
    .C(\Q[10] ),
    .D(_0294_),
    .X(_0304_));
 sky130_fd_sc_hd__and3_1 _1616_ (.A(_0880_),
    .B(sign),
    .C(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__a21oi_1 _1617_ (.A1(sign),
    .A2(_0304_),
    .B1(_0880_),
    .Y(_0306_));
 sky130_fd_sc_hd__or2_1 _1618_ (.A(net134),
    .B(net72),
    .X(_0307_));
 sky130_fd_sc_hd__o311a_1 _1619_ (.A1(_0873_),
    .A2(_0305_),
    .A3(_0306_),
    .B1(_0307_),
    .C1(_0889_),
    .X(_0140_));
 sky130_fd_sc_hd__o21ai_1 _1620_ (.A1(\Q[13] ),
    .A2(_0304_),
    .B1(sign),
    .Y(_0308_));
 sky130_fd_sc_hd__xnor2_1 _1621_ (.A(\Q[14] ),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__or2_1 _1622_ (.A(net135),
    .B(net73),
    .X(_0310_));
 sky130_fd_sc_hd__o211a_1 _1623_ (.A1(_0873_),
    .A2(_0309_),
    .B1(_0310_),
    .C1(_0889_),
    .X(_0141_));
 sky130_fd_sc_hd__o31a_1 _1624_ (.A1(\Q[14] ),
    .A2(\Q[13] ),
    .A3(_0304_),
    .B1(sign),
    .X(_0311_));
 sky130_fd_sc_hd__xor2_1 _1625_ (.A(\Q[15] ),
    .B(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__or2_1 _1626_ (.A(net134),
    .B(net74),
    .X(_0313_));
 sky130_fd_sc_hd__o211a_1 _1627_ (.A1(_0873_),
    .A2(_0312_),
    .B1(_0313_),
    .C1(_0889_),
    .X(_0142_));
 sky130_fd_sc_hd__or4_4 _1628_ (.A(\Q[15] ),
    .B(\Q[14] ),
    .C(\Q[13] ),
    .D(_0304_),
    .X(_0314_));
 sky130_fd_sc_hd__and3_1 _1629_ (.A(\Q[16] ),
    .B(sign),
    .C(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__a21oi_1 _1630_ (.A1(sign),
    .A2(_0314_),
    .B1(\Q[16] ),
    .Y(_0316_));
 sky130_fd_sc_hd__o21ai_1 _1631_ (.A1(_0315_),
    .A2(_0316_),
    .B1(net134),
    .Y(_0317_));
 sky130_fd_sc_hd__o211a_1 _1632_ (.A1(net134),
    .A2(net75),
    .B1(_0889_),
    .C1(_0317_),
    .X(_0143_));
 sky130_fd_sc_hd__o21ai_1 _1633_ (.A1(\Q[16] ),
    .A2(_0314_),
    .B1(sign),
    .Y(_0318_));
 sky130_fd_sc_hd__xnor2_1 _1634_ (.A(\Q[17] ),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__or2_1 _1635_ (.A(net134),
    .B(net76),
    .X(_0320_));
 sky130_fd_sc_hd__o211a_1 _1636_ (.A1(_0873_),
    .A2(_0319_),
    .B1(_0320_),
    .C1(_0889_),
    .X(_0144_));
 sky130_fd_sc_hd__or3_1 _1637_ (.A(\Q[17] ),
    .B(\Q[16] ),
    .C(_0314_),
    .X(_0321_));
 sky130_fd_sc_hd__nand2_1 _1638_ (.A(sign),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__and2_1 _1639_ (.A(\Q[18] ),
    .B(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__o21ai_1 _1640_ (.A1(\Q[18] ),
    .A2(_0322_),
    .B1(net134),
    .Y(_0324_));
 sky130_fd_sc_hd__o221a_1 _1641_ (.A1(net134),
    .A2(net77),
    .B1(_0323_),
    .B2(_0324_),
    .C1(_0889_),
    .X(_0145_));
 sky130_fd_sc_hd__o21ai_1 _1642_ (.A1(\Q[18] ),
    .A2(_0321_),
    .B1(sign),
    .Y(_0325_));
 sky130_fd_sc_hd__xnor2_1 _1643_ (.A(\Q[19] ),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__or2_1 _1644_ (.A(net134),
    .B(net78),
    .X(_0327_));
 sky130_fd_sc_hd__o211a_1 _1645_ (.A1(_0873_),
    .A2(_0326_),
    .B1(_0327_),
    .C1(_0889_),
    .X(_0146_));
 sky130_fd_sc_hd__o31a_1 _1646_ (.A1(\Q[19] ),
    .A2(\Q[18] ),
    .A3(_0321_),
    .B1(sign),
    .X(_0328_));
 sky130_fd_sc_hd__xor2_1 _1647_ (.A(\Q[20] ),
    .B(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__or2_1 _1648_ (.A(net134),
    .B(net80),
    .X(_0330_));
 sky130_fd_sc_hd__o211a_1 _1649_ (.A1(_0873_),
    .A2(_0329_),
    .B1(_0330_),
    .C1(_0889_),
    .X(_0147_));
 sky130_fd_sc_hd__a21oi_1 _1650_ (.A1(\Q[20] ),
    .A2(sign),
    .B1(_0328_),
    .Y(_0331_));
 sky130_fd_sc_hd__nor2_1 _1651_ (.A(\Q[21] ),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__a21o_1 _1652_ (.A1(\Q[21] ),
    .A2(_0331_),
    .B1(_0873_),
    .X(_0333_));
 sky130_fd_sc_hd__o221a_1 _1653_ (.A1(net134),
    .A2(net81),
    .B1(_0332_),
    .B2(_0333_),
    .C1(_0889_),
    .X(_0148_));
 sky130_fd_sc_hd__or4_1 _1654_ (.A(\Q[21] ),
    .B(\Q[20] ),
    .C(\Q[19] ),
    .D(\Q[18] ),
    .X(_0334_));
 sky130_fd_sc_hd__or2_1 _1655_ (.A(_0321_),
    .B(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__a21oi_1 _1656_ (.A1(sign),
    .A2(_0335_),
    .B1(_0879_),
    .Y(_0336_));
 sky130_fd_sc_hd__a31o_1 _1657_ (.A1(_0879_),
    .A2(sign),
    .A3(_0335_),
    .B1(_0873_),
    .X(_0337_));
 sky130_fd_sc_hd__o221a_1 _1658_ (.A1(net134),
    .A2(net82),
    .B1(_0336_),
    .B2(_0337_),
    .C1(_0889_),
    .X(_0149_));
 sky130_fd_sc_hd__or3_1 _1659_ (.A(\Q[22] ),
    .B(\Q[17] ),
    .C(_0334_),
    .X(_0338_));
 sky130_fd_sc_hd__o31a_1 _1660_ (.A1(\Q[16] ),
    .A2(_0314_),
    .A3(_0338_),
    .B1(sign),
    .X(_0339_));
 sky130_fd_sc_hd__xor2_1 _1661_ (.A(\Q[23] ),
    .B(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _1662_ (.A(net134),
    .B(net83),
    .X(_0341_));
 sky130_fd_sc_hd__o211a_1 _1663_ (.A1(_0873_),
    .A2(_0340_),
    .B1(_0341_),
    .C1(_0889_),
    .X(_0150_));
 sky130_fd_sc_hd__or3_1 _1664_ (.A(\Q[23] ),
    .B(\Q[16] ),
    .C(_0338_),
    .X(_0342_));
 sky130_fd_sc_hd__or2_2 _1665_ (.A(_0314_),
    .B(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__a21oi_1 _1666_ (.A1(sign),
    .A2(_0343_),
    .B1(_0878_),
    .Y(_0344_));
 sky130_fd_sc_hd__a31o_1 _1667_ (.A1(_0878_),
    .A2(sign),
    .A3(_0343_),
    .B1(_0873_),
    .X(_0345_));
 sky130_fd_sc_hd__o221a_1 _1668_ (.A1(net134),
    .A2(net84),
    .B1(_0344_),
    .B2(_0345_),
    .C1(_0889_),
    .X(_0151_));
 sky130_fd_sc_hd__o21ai_1 _1669_ (.A1(\Q[24] ),
    .A2(_0343_),
    .B1(sign),
    .Y(_0346_));
 sky130_fd_sc_hd__xnor2_1 _1670_ (.A(\Q[25] ),
    .B(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__or2_1 _1671_ (.A(net134),
    .B(net85),
    .X(_0348_));
 sky130_fd_sc_hd__o211a_1 _1672_ (.A1(_0873_),
    .A2(_0347_),
    .B1(_0348_),
    .C1(_0889_),
    .X(_0152_));
 sky130_fd_sc_hd__o31a_1 _1673_ (.A1(\Q[25] ),
    .A2(\Q[24] ),
    .A3(_0343_),
    .B1(sign),
    .X(_0349_));
 sky130_fd_sc_hd__xor2_1 _1674_ (.A(\Q[26] ),
    .B(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__or2_1 _1675_ (.A(net134),
    .B(net86),
    .X(_0351_));
 sky130_fd_sc_hd__o211a_1 _1676_ (.A1(_0873_),
    .A2(_0350_),
    .B1(_0351_),
    .C1(_0889_),
    .X(_0153_));
 sky130_fd_sc_hd__o41a_1 _1677_ (.A1(\Q[26] ),
    .A2(\Q[25] ),
    .A3(\Q[24] ),
    .A4(_0343_),
    .B1(sign),
    .X(_0352_));
 sky130_fd_sc_hd__xor2_1 _1678_ (.A(\Q[27] ),
    .B(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__or2_1 _1679_ (.A(net134),
    .B(net87),
    .X(_0354_));
 sky130_fd_sc_hd__o211a_1 _1680_ (.A1(_0873_),
    .A2(_0353_),
    .B1(_0354_),
    .C1(_0889_),
    .X(_0154_));
 sky130_fd_sc_hd__or4_1 _1681_ (.A(\Q[27] ),
    .B(\Q[26] ),
    .C(\Q[25] ),
    .D(\Q[24] ),
    .X(_0355_));
 sky130_fd_sc_hd__or2_2 _1682_ (.A(_0343_),
    .B(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__a21oi_1 _1683_ (.A1(sign),
    .A2(_0356_),
    .B1(_0877_),
    .Y(_0357_));
 sky130_fd_sc_hd__a31o_1 _1684_ (.A1(_0877_),
    .A2(sign),
    .A3(_0356_),
    .B1(_0873_),
    .X(_0358_));
 sky130_fd_sc_hd__o221a_1 _1685_ (.A1(net134),
    .A2(net88),
    .B1(_0357_),
    .B2(_0358_),
    .C1(_0889_),
    .X(_0155_));
 sky130_fd_sc_hd__o21ai_1 _1686_ (.A1(\Q[28] ),
    .A2(_0356_),
    .B1(sign),
    .Y(_0359_));
 sky130_fd_sc_hd__nor2_1 _1687_ (.A(\Q[29] ),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__a21o_1 _1688_ (.A1(\Q[29] ),
    .A2(_0359_),
    .B1(_0873_),
    .X(_0361_));
 sky130_fd_sc_hd__o221a_1 _1689_ (.A1(net135),
    .A2(net89),
    .B1(_0360_),
    .B2(_0361_),
    .C1(_0889_),
    .X(_0156_));
 sky130_fd_sc_hd__o31a_1 _1690_ (.A1(\Q[29] ),
    .A2(\Q[28] ),
    .A3(_0356_),
    .B1(sign),
    .X(_0362_));
 sky130_fd_sc_hd__xor2_1 _1691_ (.A(\Q[30] ),
    .B(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__or2_1 _1692_ (.A(net135),
    .B(net91),
    .X(_0364_));
 sky130_fd_sc_hd__o211a_1 _1693_ (.A1(_0873_),
    .A2(_0363_),
    .B1(_0364_),
    .C1(_0889_),
    .X(_0157_));
 sky130_fd_sc_hd__o41a_1 _1694_ (.A1(\Q[30] ),
    .A2(\Q[29] ),
    .A3(\Q[28] ),
    .A4(_0356_),
    .B1(sign),
    .X(_0365_));
 sky130_fd_sc_hd__xor2_1 _1695_ (.A(\Q[31] ),
    .B(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__or2_1 _1696_ (.A(net135),
    .B(net92),
    .X(_0367_));
 sky130_fd_sc_hd__o211a_1 _1697_ (.A1(_0873_),
    .A2(_0366_),
    .B1(_0367_),
    .C1(_0889_),
    .X(_0158_));
 sky130_fd_sc_hd__or4_1 _1698_ (.A(\Q[31] ),
    .B(\Q[30] ),
    .C(\Q[29] ),
    .D(\Q[28] ),
    .X(_0368_));
 sky130_fd_sc_hd__or4_2 _1699_ (.A(_0314_),
    .B(_0342_),
    .C(_0355_),
    .D(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__nand2_1 _1700_ (.A(sign),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__or3_1 _1701_ (.A(\A[0] ),
    .B(_0873_),
    .C(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__and3_1 _1702_ (.A(\A[0] ),
    .B(\count[5] ),
    .C(_0370_),
    .X(_0372_));
 sky130_fd_sc_hd__a21oi_1 _1703_ (.A1(_0873_),
    .A2(net93),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__a21oi_1 _1704_ (.A1(_0371_),
    .A2(_0373_),
    .B1(net66),
    .Y(_0159_));
 sky130_fd_sc_hd__or2_1 _1705_ (.A(\A[0] ),
    .B(_0369_),
    .X(_0374_));
 sky130_fd_sc_hd__nand2_1 _1706_ (.A(sign),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__or3_1 _1707_ (.A(\A[1] ),
    .B(_0873_),
    .C(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__and3_1 _1708_ (.A(\A[1] ),
    .B(\count[5] ),
    .C(_0375_),
    .X(_0377_));
 sky130_fd_sc_hd__a21oi_1 _1709_ (.A1(_0873_),
    .A2(net94),
    .B1(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__a21oi_1 _1710_ (.A1(_0376_),
    .A2(_0378_),
    .B1(net66),
    .Y(_0160_));
 sky130_fd_sc_hd__or2_1 _1711_ (.A(\A[1] ),
    .B(_0374_),
    .X(_0379_));
 sky130_fd_sc_hd__a21oi_1 _1712_ (.A1(sign),
    .A2(_0379_),
    .B1(_0873_),
    .Y(_0380_));
 sky130_fd_sc_hd__and4b_1 _1713_ (.A_N(\A[2] ),
    .B(net135),
    .C(sign),
    .D(_0379_),
    .X(_0381_));
 sky130_fd_sc_hd__a22o_1 _1714_ (.A1(_0873_),
    .A2(net95),
    .B1(_0380_),
    .B2(\A[2] ),
    .X(_0382_));
 sky130_fd_sc_hd__o21a_1 _1715_ (.A1(_0381_),
    .A2(_0382_),
    .B1(_0889_),
    .X(_0161_));
 sky130_fd_sc_hd__o21ai_1 _1716_ (.A1(\A[2] ),
    .A2(_0379_),
    .B1(sign),
    .Y(_0383_));
 sky130_fd_sc_hd__and3_1 _1717_ (.A(\A[3] ),
    .B(net135),
    .C(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__or3_1 _1718_ (.A(\A[3] ),
    .B(_0873_),
    .C(_0383_),
    .X(_0385_));
 sky130_fd_sc_hd__a21oi_1 _1719_ (.A1(_0873_),
    .A2(net96),
    .B1(_0384_),
    .Y(_0386_));
 sky130_fd_sc_hd__a21oi_1 _1720_ (.A1(_0385_),
    .A2(_0386_),
    .B1(net66),
    .Y(_0162_));
 sky130_fd_sc_hd__o31a_1 _1721_ (.A1(\A[3] ),
    .A2(\A[2] ),
    .A3(_0379_),
    .B1(sign),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_1 _1722_ (.A(\A[4] ),
    .B(net135),
    .Y(_0388_));
 sky130_fd_sc_hd__or3b_1 _1723_ (.A(\A[4] ),
    .B(_0873_),
    .C_N(_0387_),
    .X(_0389_));
 sky130_fd_sc_hd__o2bb2a_1 _1724_ (.A1_N(_0873_),
    .A2_N(net97),
    .B1(_0387_),
    .B2(_0388_),
    .X(_0390_));
 sky130_fd_sc_hd__a21oi_1 _1725_ (.A1(_0389_),
    .A2(_0390_),
    .B1(net66),
    .Y(_0163_));
 sky130_fd_sc_hd__a21oi_1 _1726_ (.A1(\A[4] ),
    .A2(sign),
    .B1(_0387_),
    .Y(_0391_));
 sky130_fd_sc_hd__and3_1 _1727_ (.A(\A[5] ),
    .B(net135),
    .C(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__or2_1 _1728_ (.A(\A[5] ),
    .B(_0873_),
    .X(_0393_));
 sky130_fd_sc_hd__a2bb2o_1 _1729_ (.A1_N(_0393_),
    .A2_N(_0391_),
    .B1(net98),
    .B2(_0873_),
    .X(_0394_));
 sky130_fd_sc_hd__o21a_1 _1730_ (.A1(_0392_),
    .A2(_0394_),
    .B1(_0889_),
    .X(_0164_));
 sky130_fd_sc_hd__or4_1 _1731_ (.A(\A[5] ),
    .B(\A[4] ),
    .C(\A[3] ),
    .D(\A[2] ),
    .X(_0395_));
 sky130_fd_sc_hd__o21a_1 _1732_ (.A1(_0379_),
    .A2(_0395_),
    .B1(sign),
    .X(_0396_));
 sky130_fd_sc_hd__nand2_1 _1733_ (.A(\count[5] ),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__or3b_1 _1734_ (.A(_0396_),
    .B(_0873_),
    .C_N(\A[6] ),
    .X(_0398_));
 sky130_fd_sc_hd__o221a_1 _1735_ (.A1(\count[5] ),
    .A2(_0876_),
    .B1(_0397_),
    .B2(\A[6] ),
    .C1(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__nor2_1 _1736_ (.A(net66),
    .B(_0399_),
    .Y(_0165_));
 sky130_fd_sc_hd__or4_1 _1737_ (.A(\A[6] ),
    .B(\A[1] ),
    .C(_0374_),
    .D(_0395_),
    .X(_0400_));
 sky130_fd_sc_hd__a21oi_1 _1738_ (.A1(sign),
    .A2(_0400_),
    .B1(_0873_),
    .Y(_0401_));
 sky130_fd_sc_hd__and4b_1 _1739_ (.A_N(\A[7] ),
    .B(\count[5] ),
    .C(sign),
    .D(_0400_),
    .X(_0402_));
 sky130_fd_sc_hd__a22o_1 _1740_ (.A1(_0873_),
    .A2(net100),
    .B1(_0401_),
    .B2(\A[7] ),
    .X(_0403_));
 sky130_fd_sc_hd__o21a_1 _1741_ (.A1(_0402_),
    .A2(_0403_),
    .B1(_0889_),
    .X(_0166_));
 sky130_fd_sc_hd__or2_1 _1742_ (.A(\A[7] ),
    .B(\A[0] ),
    .X(_0404_));
 sky130_fd_sc_hd__or4_1 _1743_ (.A(\A[6] ),
    .B(\A[1] ),
    .C(_0395_),
    .D(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__or2_1 _1744_ (.A(_0369_),
    .B(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__nand2_1 _1745_ (.A(sign),
    .B(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__nor3_1 _1746_ (.A(\A[8] ),
    .B(_0873_),
    .C(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__and2_1 _1747_ (.A(_0873_),
    .B(net102),
    .X(_0409_));
 sky130_fd_sc_hd__a31o_1 _1748_ (.A1(\A[8] ),
    .A2(\count[5] ),
    .A3(_0407_),
    .B1(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__o21a_1 _1749_ (.A1(_0408_),
    .A2(_0410_),
    .B1(_0889_),
    .X(_0167_));
 sky130_fd_sc_hd__o21ai_1 _1750_ (.A1(\A[8] ),
    .A2(_0406_),
    .B1(sign),
    .Y(_0411_));
 sky130_fd_sc_hd__and3_1 _1751_ (.A(\A[9] ),
    .B(\count[5] ),
    .C(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__or3_1 _1752_ (.A(\A[9] ),
    .B(_0873_),
    .C(_0411_),
    .X(_0413_));
 sky130_fd_sc_hd__a21oi_1 _1753_ (.A1(_0873_),
    .A2(net103),
    .B1(_0412_),
    .Y(_0414_));
 sky130_fd_sc_hd__a21oi_1 _1754_ (.A1(_0413_),
    .A2(_0414_),
    .B1(net66),
    .Y(_0168_));
 sky130_fd_sc_hd__o31ai_1 _1755_ (.A1(\A[9] ),
    .A2(\A[8] ),
    .A3(_0406_),
    .B1(sign),
    .Y(_0415_));
 sky130_fd_sc_hd__or2_1 _1756_ (.A(\A[10] ),
    .B(_0873_),
    .X(_0416_));
 sky130_fd_sc_hd__or2_1 _1757_ (.A(_0415_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__and3_1 _1758_ (.A(\A[10] ),
    .B(\count[5] ),
    .C(_0415_),
    .X(_0418_));
 sky130_fd_sc_hd__a21oi_1 _1759_ (.A1(_0873_),
    .A2(net104),
    .B1(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__a21oi_1 _1760_ (.A1(_0417_),
    .A2(_0419_),
    .B1(net66),
    .Y(_0169_));
 sky130_fd_sc_hd__or4_1 _1761_ (.A(\A[10] ),
    .B(\A[9] ),
    .C(\A[8] ),
    .D(_0406_),
    .X(_0420_));
 sky130_fd_sc_hd__nand2_1 _1762_ (.A(sign),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__or2_1 _1763_ (.A(\A[11] ),
    .B(_0873_),
    .X(_0422_));
 sky130_fd_sc_hd__nor2_1 _1764_ (.A(_0421_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__and2_1 _1765_ (.A(_0873_),
    .B(net105),
    .X(_0424_));
 sky130_fd_sc_hd__a31o_1 _1766_ (.A1(\A[11] ),
    .A2(\count[5] ),
    .A3(_0421_),
    .B1(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__o21a_1 _1767_ (.A1(_0423_),
    .A2(_0425_),
    .B1(_0889_),
    .X(_0170_));
 sky130_fd_sc_hd__or4_1 _1768_ (.A(\A[11] ),
    .B(\A[10] ),
    .C(\A[9] ),
    .D(\A[8] ),
    .X(_0426_));
 sky130_fd_sc_hd__or3_2 _1769_ (.A(_0369_),
    .B(_0405_),
    .C(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _1770_ (.A(sign),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__or3_1 _1771_ (.A(\A[12] ),
    .B(_0873_),
    .C(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__and3_1 _1772_ (.A(\A[12] ),
    .B(\count[5] ),
    .C(_0428_),
    .X(_0430_));
 sky130_fd_sc_hd__a21oi_1 _1773_ (.A1(_0873_),
    .A2(net106),
    .B1(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__a21oi_1 _1774_ (.A1(_0429_),
    .A2(_0431_),
    .B1(net66),
    .Y(_0171_));
 sky130_fd_sc_hd__o21ai_1 _1775_ (.A1(\A[12] ),
    .A2(_0427_),
    .B1(sign),
    .Y(_0432_));
 sky130_fd_sc_hd__and3_1 _1776_ (.A(\A[13] ),
    .B(\count[5] ),
    .C(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__or3_1 _1777_ (.A(\A[13] ),
    .B(_0873_),
    .C(_0432_),
    .X(_0434_));
 sky130_fd_sc_hd__a21oi_1 _1778_ (.A1(_0873_),
    .A2(net107),
    .B1(_0433_),
    .Y(_0435_));
 sky130_fd_sc_hd__a21oi_1 _1779_ (.A1(_0434_),
    .A2(_0435_),
    .B1(net66),
    .Y(_0172_));
 sky130_fd_sc_hd__o31a_1 _1780_ (.A1(\A[13] ),
    .A2(\A[12] ),
    .A3(_0427_),
    .B1(sign),
    .X(_0436_));
 sky130_fd_sc_hd__or3b_1 _1781_ (.A(\A[14] ),
    .B(_0873_),
    .C_N(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__nand2_1 _1782_ (.A(\A[14] ),
    .B(\count[5] ),
    .Y(_0438_));
 sky130_fd_sc_hd__o2bb2a_1 _1783_ (.A1_N(_0873_),
    .A2_N(net108),
    .B1(_0436_),
    .B2(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__a21oi_1 _1784_ (.A1(_0437_),
    .A2(_0439_),
    .B1(net66),
    .Y(_0173_));
 sky130_fd_sc_hd__a21oi_1 _1785_ (.A1(\A[14] ),
    .A2(sign),
    .B1(_0436_),
    .Y(_0440_));
 sky130_fd_sc_hd__and3_1 _1786_ (.A(\A[15] ),
    .B(\count[5] ),
    .C(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__or2_1 _1787_ (.A(\A[15] ),
    .B(_0873_),
    .X(_0442_));
 sky130_fd_sc_hd__a2bb2o_1 _1788_ (.A1_N(_0442_),
    .A2_N(_0440_),
    .B1(net109),
    .B2(_0873_),
    .X(_0443_));
 sky130_fd_sc_hd__o21a_1 _1789_ (.A1(_0441_),
    .A2(_0443_),
    .B1(_0889_),
    .X(_0174_));
 sky130_fd_sc_hd__or4_1 _1790_ (.A(\A[15] ),
    .B(\A[14] ),
    .C(\A[13] ),
    .D(\A[12] ),
    .X(_0444_));
 sky130_fd_sc_hd__o21a_1 _1791_ (.A1(_0427_),
    .A2(_0444_),
    .B1(sign),
    .X(_0445_));
 sky130_fd_sc_hd__or3b_1 _1792_ (.A(\A[16] ),
    .B(_0873_),
    .C_N(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__nand2_1 _1793_ (.A(\A[16] ),
    .B(\count[5] ),
    .Y(_0447_));
 sky130_fd_sc_hd__o2bb2a_1 _1794_ (.A1_N(_0873_),
    .A2_N(net110),
    .B1(_0445_),
    .B2(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__a21oi_1 _1795_ (.A1(_0446_),
    .A2(_0448_),
    .B1(net66),
    .Y(_0175_));
 sky130_fd_sc_hd__nor3_1 _1796_ (.A(\A[16] ),
    .B(_0427_),
    .C(_0444_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2b_1 _1797_ (.A_N(_0449_),
    .B(sign),
    .Y(_0450_));
 sky130_fd_sc_hd__and3_1 _1798_ (.A(\A[17] ),
    .B(\count[5] ),
    .C(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__or3_1 _1799_ (.A(\A[17] ),
    .B(_0873_),
    .C(_0450_),
    .X(_0452_));
 sky130_fd_sc_hd__a21oi_1 _1800_ (.A1(_0873_),
    .A2(net111),
    .B1(_0451_),
    .Y(_0453_));
 sky130_fd_sc_hd__a21oi_1 _1801_ (.A1(_0452_),
    .A2(_0453_),
    .B1(net66),
    .Y(_0176_));
 sky130_fd_sc_hd__o41a_1 _1802_ (.A1(\A[17] ),
    .A2(\A[16] ),
    .A3(_0427_),
    .A4(_0444_),
    .B1(sign),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_1 _1803_ (.A(\A[18] ),
    .B(net134),
    .Y(_0455_));
 sky130_fd_sc_hd__or3b_1 _1804_ (.A(\A[18] ),
    .B(_0873_),
    .C_N(_0454_),
    .X(_0456_));
 sky130_fd_sc_hd__o2bb2a_1 _1805_ (.A1_N(_0873_),
    .A2_N(net113),
    .B1(_0454_),
    .B2(_0455_),
    .X(_0457_));
 sky130_fd_sc_hd__a21oi_1 _1806_ (.A1(_0456_),
    .A2(_0457_),
    .B1(net66),
    .Y(_0177_));
 sky130_fd_sc_hd__a21oi_1 _1807_ (.A1(\A[18] ),
    .A2(sign),
    .B1(_0454_),
    .Y(_0458_));
 sky130_fd_sc_hd__and3_1 _1808_ (.A(\A[19] ),
    .B(net134),
    .C(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__or3_1 _1809_ (.A(\A[19] ),
    .B(_0873_),
    .C(_0458_),
    .X(_0460_));
 sky130_fd_sc_hd__a21oi_1 _1810_ (.A1(_0873_),
    .A2(net114),
    .B1(_0459_),
    .Y(_0461_));
 sky130_fd_sc_hd__a21oi_1 _1811_ (.A1(_0460_),
    .A2(_0461_),
    .B1(net66),
    .Y(_0178_));
 sky130_fd_sc_hd__or2_1 _1812_ (.A(\A[19] ),
    .B(\A[18] ),
    .X(_0462_));
 sky130_fd_sc_hd__a21o_1 _1813_ (.A1(sign),
    .A2(_0462_),
    .B1(_0454_),
    .X(_0463_));
 sky130_fd_sc_hd__nand2_1 _1814_ (.A(\A[20] ),
    .B(net134),
    .Y(_0464_));
 sky130_fd_sc_hd__or3b_1 _1815_ (.A(\A[20] ),
    .B(_0873_),
    .C_N(_0463_),
    .X(_0465_));
 sky130_fd_sc_hd__o2bb2a_1 _1816_ (.A1_N(_0873_),
    .A2_N(net115),
    .B1(_0463_),
    .B2(_0464_),
    .X(_0466_));
 sky130_fd_sc_hd__a21oi_1 _1817_ (.A1(_0465_),
    .A2(_0466_),
    .B1(net66),
    .Y(_0179_));
 sky130_fd_sc_hd__a21oi_1 _1818_ (.A1(\A[20] ),
    .A2(sign),
    .B1(_0463_),
    .Y(_0467_));
 sky130_fd_sc_hd__nand3_1 _1819_ (.A(\A[21] ),
    .B(net134),
    .C(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_1 _1820_ (.A(_0873_),
    .B(net116),
    .Y(_0469_));
 sky130_fd_sc_hd__o311a_1 _1821_ (.A1(\A[21] ),
    .A2(_0873_),
    .A3(_0467_),
    .B1(_0468_),
    .C1(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__nor2_1 _1822_ (.A(net66),
    .B(_0470_),
    .Y(_0180_));
 sky130_fd_sc_hd__or3_1 _1823_ (.A(\A[21] ),
    .B(\A[20] ),
    .C(_0462_),
    .X(_0471_));
 sky130_fd_sc_hd__a21o_1 _1824_ (.A1(sign),
    .A2(_0471_),
    .B1(_0454_),
    .X(_0472_));
 sky130_fd_sc_hd__nand2_1 _1825_ (.A(\A[22] ),
    .B(net134),
    .Y(_0473_));
 sky130_fd_sc_hd__or3b_1 _1826_ (.A(\A[22] ),
    .B(_0873_),
    .C_N(_0472_),
    .X(_0474_));
 sky130_fd_sc_hd__o221a_1 _1827_ (.A1(net134),
    .A2(_0875_),
    .B1(_0472_),
    .B2(_0473_),
    .C1(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__nor2_1 _1828_ (.A(net66),
    .B(_0475_),
    .Y(_0181_));
 sky130_fd_sc_hd__or2_1 _1829_ (.A(\A[22] ),
    .B(_0471_),
    .X(_0476_));
 sky130_fd_sc_hd__a21oi_1 _1830_ (.A1(\A[22] ),
    .A2(sign),
    .B1(_0472_),
    .Y(_0477_));
 sky130_fd_sc_hd__or3_1 _1831_ (.A(\A[23] ),
    .B(_0873_),
    .C(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__and3_1 _1832_ (.A(\A[23] ),
    .B(net134),
    .C(_0477_),
    .X(_0479_));
 sky130_fd_sc_hd__a21oi_1 _1833_ (.A1(_0873_),
    .A2(net118),
    .B1(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a21oi_1 _1834_ (.A1(_0478_),
    .A2(_0480_),
    .B1(net66),
    .Y(_0182_));
 sky130_fd_sc_hd__or4b_2 _1835_ (.A(\A[23] ),
    .B(_0476_),
    .C(\A[17] ),
    .D_N(_0449_),
    .X(_0481_));
 sky130_fd_sc_hd__nand2_1 _1836_ (.A(sign),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__or2_1 _1837_ (.A(\A[24] ),
    .B(_0873_),
    .X(_0483_));
 sky130_fd_sc_hd__a2bb2o_1 _1838_ (.A1_N(_0482_),
    .A2_N(_0483_),
    .B1(_0873_),
    .B2(net119),
    .X(_0484_));
 sky130_fd_sc_hd__a31o_1 _1839_ (.A1(\A[24] ),
    .A2(net134),
    .A3(_0482_),
    .B1(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__and2_1 _1840_ (.A(_0889_),
    .B(_0485_),
    .X(_0183_));
 sky130_fd_sc_hd__o21ai_1 _1841_ (.A1(\A[24] ),
    .A2(_0481_),
    .B1(sign),
    .Y(_0486_));
 sky130_fd_sc_hd__and3_1 _1842_ (.A(\A[25] ),
    .B(net134),
    .C(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__or3_1 _1843_ (.A(\A[25] ),
    .B(_0873_),
    .C(_0486_),
    .X(_0488_));
 sky130_fd_sc_hd__a21oi_1 _1844_ (.A1(_0873_),
    .A2(net120),
    .B1(_0487_),
    .Y(_0489_));
 sky130_fd_sc_hd__a21oi_1 _1845_ (.A1(_0488_),
    .A2(_0489_),
    .B1(net66),
    .Y(_0184_));
 sky130_fd_sc_hd__o31a_1 _1846_ (.A1(\A[25] ),
    .A2(\A[24] ),
    .A3(_0481_),
    .B1(sign),
    .X(_0490_));
 sky130_fd_sc_hd__or3b_1 _1847_ (.A(\A[26] ),
    .B(_0873_),
    .C_N(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__nand2_1 _1848_ (.A(\A[26] ),
    .B(net134),
    .Y(_0492_));
 sky130_fd_sc_hd__o2bb2a_1 _1849_ (.A1_N(_0873_),
    .A2_N(net121),
    .B1(_0490_),
    .B2(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__a21oi_1 _1850_ (.A1(_0491_),
    .A2(_0493_),
    .B1(net66),
    .Y(_0185_));
 sky130_fd_sc_hd__a21oi_1 _1851_ (.A1(\A[26] ),
    .A2(sign),
    .B1(_0490_),
    .Y(_0494_));
 sky130_fd_sc_hd__and3_1 _1852_ (.A(\A[27] ),
    .B(net134),
    .C(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__or3_1 _1853_ (.A(\A[27] ),
    .B(_0873_),
    .C(_0494_),
    .X(_0496_));
 sky130_fd_sc_hd__a21oi_1 _1854_ (.A1(_0873_),
    .A2(net122),
    .B1(_0495_),
    .Y(_0497_));
 sky130_fd_sc_hd__a21oi_1 _1855_ (.A1(_0496_),
    .A2(_0497_),
    .B1(net66),
    .Y(_0186_));
 sky130_fd_sc_hd__or4_1 _1856_ (.A(\A[27] ),
    .B(\A[26] ),
    .C(\A[25] ),
    .D(\A[24] ),
    .X(_0498_));
 sky130_fd_sc_hd__o21a_1 _1857_ (.A1(_0481_),
    .A2(_0498_),
    .B1(sign),
    .X(_0499_));
 sky130_fd_sc_hd__or3b_1 _1858_ (.A(\A[28] ),
    .B(_0873_),
    .C_N(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__nand2_1 _1859_ (.A(\A[28] ),
    .B(net134),
    .Y(_0501_));
 sky130_fd_sc_hd__o2bb2a_1 _1860_ (.A1_N(_0873_),
    .A2_N(net124),
    .B1(_0499_),
    .B2(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__a21oi_1 _1861_ (.A1(_0500_),
    .A2(_0502_),
    .B1(net66),
    .Y(_0187_));
 sky130_fd_sc_hd__a21oi_1 _1862_ (.A1(\A[28] ),
    .A2(sign),
    .B1(_0499_),
    .Y(_0503_));
 sky130_fd_sc_hd__and3_1 _1863_ (.A(\A[29] ),
    .B(net134),
    .C(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__or3_1 _1864_ (.A(\A[29] ),
    .B(_0873_),
    .C(_0503_),
    .X(_0505_));
 sky130_fd_sc_hd__a21oi_1 _1865_ (.A1(_0873_),
    .A2(net125),
    .B1(_0504_),
    .Y(_0506_));
 sky130_fd_sc_hd__a21oi_1 _1866_ (.A1(_0505_),
    .A2(_0506_),
    .B1(net66),
    .Y(_0188_));
 sky130_fd_sc_hd__or4_1 _1867_ (.A(\A[29] ),
    .B(\A[28] ),
    .C(_0481_),
    .D(_0498_),
    .X(_0507_));
 sky130_fd_sc_hd__nand2_1 _1868_ (.A(sign),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__or3_1 _1869_ (.A(\A[30] ),
    .B(_0873_),
    .C(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__and3_1 _1870_ (.A(\A[30] ),
    .B(net134),
    .C(_0508_),
    .X(_0510_));
 sky130_fd_sc_hd__a21oi_1 _1871_ (.A1(_0873_),
    .A2(net126),
    .B1(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__a21oi_1 _1872_ (.A1(_0509_),
    .A2(_0511_),
    .B1(net66),
    .Y(_0189_));
 sky130_fd_sc_hd__a21boi_1 _1873_ (.A1(\A[30] ),
    .A2(sign),
    .B1_N(_0508_),
    .Y(_0512_));
 sky130_fd_sc_hd__nand3_1 _1874_ (.A(\A[31] ),
    .B(net134),
    .C(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_1 _1875_ (.A(_0873_),
    .B(net127),
    .Y(_0514_));
 sky130_fd_sc_hd__o311a_1 _1876_ (.A1(\A[31] ),
    .A2(_0873_),
    .A3(_0512_),
    .B1(_0513_),
    .C1(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__nor2_1 _1877_ (.A(net66),
    .B(_0515_),
    .Y(_0190_));
 sky130_fd_sc_hd__o21a_1 _1878_ (.A1(net135),
    .A2(net67),
    .B1(_0889_),
    .X(_0191_));
 sky130_fd_sc_hd__o32a_1 _1879_ (.A1(net25),
    .A2(_0891_),
    .A3(_1044_),
    .B1(_0888_),
    .B2(net66),
    .X(_0516_));
 sky130_fd_sc_hd__inv_2 _1880_ (.A(_0516_),
    .Y(_0192_));
 sky130_fd_sc_hd__or4_1 _1881_ (.A(net55),
    .B(net57),
    .C(_0890_),
    .D(_0966_),
    .X(_0517_));
 sky130_fd_sc_hd__a21bo_1 _1882_ (.A1(\abs_multiplier[31] ),
    .A2(_0889_),
    .B1_N(_0517_),
    .X(_0193_));
 sky130_fd_sc_hd__a21oi_1 _1883_ (.A1(_0873_),
    .A2(\count[0] ),
    .B1(net66),
    .Y(_0518_));
 sky130_fd_sc_hd__o21a_1 _1884_ (.A1(_0873_),
    .A2(\count[0] ),
    .B1(_0518_),
    .X(_0194_));
 sky130_fd_sc_hd__a21oi_1 _1885_ (.A1(_0873_),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .Y(_0519_));
 sky130_fd_sc_hd__and3_1 _1886_ (.A(_0873_),
    .B(\count[1] ),
    .C(\count[0] ),
    .X(_0520_));
 sky130_fd_sc_hd__nor3_1 _1887_ (.A(net66),
    .B(_0519_),
    .C(_0520_),
    .Y(_0195_));
 sky130_fd_sc_hd__and2_1 _1888_ (.A(\count[2] ),
    .B(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__nor2_1 _1889_ (.A(net66),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__o21a_1 _1890_ (.A1(\count[2] ),
    .A2(_0520_),
    .B1(_0522_),
    .X(_0196_));
 sky130_fd_sc_hd__and3_1 _1891_ (.A(\count[3] ),
    .B(\count[2] ),
    .C(_0520_),
    .X(_0523_));
 sky130_fd_sc_hd__nor2_1 _1892_ (.A(net66),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__o21a_1 _1893_ (.A1(\count[3] ),
    .A2(_0521_),
    .B1(_0524_),
    .X(_0197_));
 sky130_fd_sc_hd__a21oi_1 _1894_ (.A1(\count[4] ),
    .A2(_0523_),
    .B1(net66),
    .Y(_0525_));
 sky130_fd_sc_hd__o21a_1 _1895_ (.A1(\count[4] ),
    .A2(_0523_),
    .B1(_0525_),
    .X(_0198_));
 sky130_fd_sc_hd__a41o_1 _1896_ (.A1(\count[3] ),
    .A2(\count[2] ),
    .A3(\count[1] ),
    .A4(\count[0] ),
    .B1(net135),
    .X(_0526_));
 sky130_fd_sc_hd__and3_1 _1897_ (.A(_0889_),
    .B(_1047_),
    .C(_0526_),
    .X(_0199_));
 sky130_fd_sc_hd__nor2_1 _1898_ (.A(\A[1] ),
    .B(_1054_),
    .Y(_0527_));
 sky130_fd_sc_hd__o211ai_1 _1899_ (.A1(_0883_),
    .A2(_1049_),
    .B1(_1052_),
    .C1(_0872_),
    .Y(_0528_));
 sky130_fd_sc_hd__o211a_1 _1900_ (.A1(\M[1] ),
    .A2(_1049_),
    .B1(_1053_),
    .C1(\A[1] ),
    .X(_0529_));
 sky130_fd_sc_hd__nor2_1 _1901_ (.A(_0527_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__and2_1 _1902_ (.A(\A[0] ),
    .B(_1051_),
    .X(_0531_));
 sky130_fd_sc_hd__nand2_1 _1903_ (.A(_0530_),
    .B(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__o21a_1 _1904_ (.A1(_0530_),
    .A2(_0531_),
    .B1(_1148_),
    .X(_0533_));
 sky130_fd_sc_hd__a221o_1 _1905_ (.A1(\A[1] ),
    .A2(_1149_),
    .B1(_0532_),
    .B2(_0533_),
    .C1(\count[5] ),
    .X(_0534_));
 sky130_fd_sc_hd__o211a_1 _1906_ (.A1(\A[0] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0534_),
    .X(_0200_));
 sky130_fd_sc_hd__a31o_1 _1907_ (.A1(\A[0] ),
    .A2(_1051_),
    .A3(_0528_),
    .B1(_0529_),
    .X(_0535_));
 sky130_fd_sc_hd__xor2_1 _1908_ (.A(\A[2] ),
    .B(_1055_),
    .X(_0536_));
 sky130_fd_sc_hd__nand2_1 _1909_ (.A(_0535_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__o21a_1 _1910_ (.A1(_0535_),
    .A2(_0536_),
    .B1(_1148_),
    .X(_0538_));
 sky130_fd_sc_hd__a221o_1 _1911_ (.A1(\A[2] ),
    .A2(_1149_),
    .B1(_0537_),
    .B2(_0538_),
    .C1(net135),
    .X(_0539_));
 sky130_fd_sc_hd__o211a_1 _1912_ (.A1(\A[1] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0539_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_1 _1913_ (.A(\A[3] ),
    .B(_1056_),
    .X(_0540_));
 sky130_fd_sc_hd__xor2_1 _1914_ (.A(\A[3] ),
    .B(_1056_),
    .X(_0541_));
 sky130_fd_sc_hd__a21bo_1 _1915_ (.A1(\A[2] ),
    .A2(_1055_),
    .B1_N(_0537_),
    .X(_0542_));
 sky130_fd_sc_hd__a21oi_1 _1916_ (.A1(_0541_),
    .A2(_0542_),
    .B1(_1149_),
    .Y(_0543_));
 sky130_fd_sc_hd__o21a_1 _1917_ (.A1(_0541_),
    .A2(_0542_),
    .B1(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__a21o_1 _1918_ (.A1(\A[3] ),
    .A2(_1149_),
    .B1(net135),
    .X(_0545_));
 sky130_fd_sc_hd__o221a_1 _1919_ (.A1(\A[2] ),
    .A2(_0873_),
    .B1(_0544_),
    .B2(_0545_),
    .C1(_0889_),
    .X(_0202_));
 sky130_fd_sc_hd__xor2_1 _1920_ (.A(\A[4] ),
    .B(_1057_),
    .X(_0546_));
 sky130_fd_sc_hd__o211a_1 _1921_ (.A1(\A[3] ),
    .A2(_1056_),
    .B1(_1055_),
    .C1(\A[2] ),
    .X(_0547_));
 sky130_fd_sc_hd__a311o_1 _1922_ (.A1(_0535_),
    .A2(_0536_),
    .A3(_0541_),
    .B1(_0547_),
    .C1(_0540_),
    .X(_0548_));
 sky130_fd_sc_hd__nand2_1 _1923_ (.A(_0546_),
    .B(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__nor2_1 _1924_ (.A(_0546_),
    .B(_0548_),
    .Y(_0550_));
 sky130_fd_sc_hd__and3b_1 _1925_ (.A_N(_0550_),
    .B(_1148_),
    .C(_0549_),
    .X(_0551_));
 sky130_fd_sc_hd__a21o_1 _1926_ (.A1(\A[4] ),
    .A2(_1149_),
    .B1(net135),
    .X(_0552_));
 sky130_fd_sc_hd__o221a_1 _1927_ (.A1(\A[3] ),
    .A2(_0873_),
    .B1(_0551_),
    .B2(_0552_),
    .C1(_0889_),
    .X(_0203_));
 sky130_fd_sc_hd__nor2_1 _1928_ (.A(\A[5] ),
    .B(_1058_),
    .Y(_0553_));
 sky130_fd_sc_hd__xor2_1 _1929_ (.A(\A[5] ),
    .B(_1058_),
    .X(_0554_));
 sky130_fd_sc_hd__a21bo_1 _1930_ (.A1(\A[4] ),
    .A2(_1057_),
    .B1_N(_0549_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _1931_ (.A(_0554_),
    .B(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__o211a_1 _1932_ (.A1(_0554_),
    .A2(_0555_),
    .B1(_0556_),
    .C1(_1148_),
    .X(_0557_));
 sky130_fd_sc_hd__a21o_1 _1933_ (.A1(\A[5] ),
    .A2(_1149_),
    .B1(\count[5] ),
    .X(_0558_));
 sky130_fd_sc_hd__o221a_1 _1934_ (.A1(\A[4] ),
    .A2(_0873_),
    .B1(_0557_),
    .B2(_0558_),
    .C1(_0889_),
    .X(_0204_));
 sky130_fd_sc_hd__xor2_1 _1935_ (.A(\A[6] ),
    .B(_1059_),
    .X(_0559_));
 sky130_fd_sc_hd__a22oi_1 _1936_ (.A1(\A[4] ),
    .A2(_1057_),
    .B1(_1058_),
    .B2(\A[5] ),
    .Y(_0560_));
 sky130_fd_sc_hd__a21oi_1 _1937_ (.A1(_0549_),
    .A2(_0560_),
    .B1(_0553_),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_1 _1938_ (.A(_0559_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__o21a_1 _1939_ (.A1(_0559_),
    .A2(_0561_),
    .B1(_1148_),
    .X(_0563_));
 sky130_fd_sc_hd__a221o_1 _1940_ (.A1(\A[6] ),
    .A2(_1149_),
    .B1(_0562_),
    .B2(_0563_),
    .C1(\count[5] ),
    .X(_0564_));
 sky130_fd_sc_hd__and3_1 _1941_ (.A(_0889_),
    .B(_0393_),
    .C(_0564_),
    .X(_0205_));
 sky130_fd_sc_hd__xor2_1 _1942_ (.A(\A[7] ),
    .B(_1060_),
    .X(_0565_));
 sky130_fd_sc_hd__a21bo_1 _1943_ (.A1(\A[6] ),
    .A2(_1059_),
    .B1_N(_0562_),
    .X(_0566_));
 sky130_fd_sc_hd__a21oi_1 _1944_ (.A1(_0565_),
    .A2(_0566_),
    .B1(_1149_),
    .Y(_0567_));
 sky130_fd_sc_hd__o21a_1 _1945_ (.A1(_0565_),
    .A2(_0566_),
    .B1(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__a21o_1 _1946_ (.A1(\A[7] ),
    .A2(_1149_),
    .B1(\count[5] ),
    .X(_0569_));
 sky130_fd_sc_hd__o221a_1 _1947_ (.A1(\A[6] ),
    .A2(_0873_),
    .B1(_0568_),
    .B2(_0569_),
    .C1(_0889_),
    .X(_0206_));
 sky130_fd_sc_hd__and4_1 _1948_ (.A(_0546_),
    .B(_0554_),
    .C(_0559_),
    .D(_0565_),
    .X(_0570_));
 sky130_fd_sc_hd__nand2_1 _1949_ (.A(_0548_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__and4bb_1 _1950_ (.A_N(_0553_),
    .B_N(_0560_),
    .C(_0565_),
    .D(_0559_),
    .X(_0572_));
 sky130_fd_sc_hd__o211a_1 _1951_ (.A1(\A[7] ),
    .A2(_1060_),
    .B1(_1059_),
    .C1(\A[6] ),
    .X(_0573_));
 sky130_fd_sc_hd__a211oi_2 _1952_ (.A1(\A[7] ),
    .A2(_1060_),
    .B1(_0572_),
    .C1(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__xnor2_1 _1953_ (.A(\A[8] ),
    .B(_1061_),
    .Y(_0575_));
 sky130_fd_sc_hd__a21oi_1 _1954_ (.A1(_0571_),
    .A2(_0574_),
    .B1(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__a31o_1 _1955_ (.A1(_0571_),
    .A2(_0574_),
    .A3(_0575_),
    .B1(_1149_),
    .X(_0577_));
 sky130_fd_sc_hd__nor2_1 _1956_ (.A(_0576_),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__a21o_1 _1957_ (.A1(\A[8] ),
    .A2(_1149_),
    .B1(\count[5] ),
    .X(_0579_));
 sky130_fd_sc_hd__o221a_1 _1958_ (.A1(\A[7] ),
    .A2(_0873_),
    .B1(_0578_),
    .B2(_0579_),
    .C1(_0889_),
    .X(_0207_));
 sky130_fd_sc_hd__and2_1 _1959_ (.A(\A[9] ),
    .B(_1062_),
    .X(_0580_));
 sky130_fd_sc_hd__or2_1 _1960_ (.A(\A[9] ),
    .B(_1062_),
    .X(_0581_));
 sky130_fd_sc_hd__and2b_1 _1961_ (.A_N(_0580_),
    .B(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__a21o_1 _1962_ (.A1(\A[8] ),
    .A2(_1061_),
    .B1(_0576_),
    .X(_0583_));
 sky130_fd_sc_hd__a21oi_1 _1963_ (.A1(_0582_),
    .A2(_0583_),
    .B1(_1149_),
    .Y(_0584_));
 sky130_fd_sc_hd__o21a_1 _1964_ (.A1(_0582_),
    .A2(_0583_),
    .B1(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__a21o_1 _1965_ (.A1(\A[9] ),
    .A2(_1149_),
    .B1(\count[5] ),
    .X(_0586_));
 sky130_fd_sc_hd__o221a_1 _1966_ (.A1(\A[8] ),
    .A2(_0873_),
    .B1(_0585_),
    .B2(_0586_),
    .C1(_0889_),
    .X(_0208_));
 sky130_fd_sc_hd__nand2_1 _1967_ (.A(\A[10] ),
    .B(_1063_),
    .Y(_0587_));
 sky130_fd_sc_hd__xnor2_1 _1968_ (.A(\A[10] ),
    .B(_1063_),
    .Y(_0588_));
 sky130_fd_sc_hd__a21oi_1 _1969_ (.A1(_0581_),
    .A2(_0583_),
    .B1(_0580_),
    .Y(_0589_));
 sky130_fd_sc_hd__a21oi_1 _1970_ (.A1(_0588_),
    .A2(_0589_),
    .B1(_1149_),
    .Y(_0590_));
 sky130_fd_sc_hd__o21a_1 _1971_ (.A1(_0588_),
    .A2(_0589_),
    .B1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__a21o_1 _1972_ (.A1(\A[10] ),
    .A2(_1149_),
    .B1(\count[5] ),
    .X(_0592_));
 sky130_fd_sc_hd__o221a_1 _1973_ (.A1(\A[9] ),
    .A2(_0873_),
    .B1(_0591_),
    .B2(_0592_),
    .C1(_0889_),
    .X(_0209_));
 sky130_fd_sc_hd__and2_1 _1974_ (.A(\A[11] ),
    .B(_1064_),
    .X(_0593_));
 sky130_fd_sc_hd__xnor2_1 _1975_ (.A(\A[11] ),
    .B(_1064_),
    .Y(_0594_));
 sky130_fd_sc_hd__o21a_1 _1976_ (.A1(_0588_),
    .A2(_0589_),
    .B1(_0587_),
    .X(_0595_));
 sky130_fd_sc_hd__nor2_1 _1977_ (.A(_0594_),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__a21o_1 _1978_ (.A1(_0594_),
    .A2(_0595_),
    .B1(_1149_),
    .X(_0597_));
 sky130_fd_sc_hd__a2bb2o_1 _1979_ (.A1_N(_0596_),
    .A2_N(_0597_),
    .B1(\A[11] ),
    .B2(_1149_),
    .X(_0598_));
 sky130_fd_sc_hd__o211a_1 _1980_ (.A1(\count[5] ),
    .A2(_0598_),
    .B1(_0416_),
    .C1(_0889_),
    .X(_0210_));
 sky130_fd_sc_hd__and2_1 _1981_ (.A(\A[12] ),
    .B(_1065_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_1 _1982_ (.A(\A[12] ),
    .B(_1065_),
    .Y(_0600_));
 sky130_fd_sc_hd__nor2_1 _1983_ (.A(_0599_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__nor2_1 _1984_ (.A(_0588_),
    .B(_0594_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand3b_1 _1985_ (.A_N(_0575_),
    .B(_0582_),
    .C(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__a21oi_2 _1986_ (.A1(_0571_),
    .A2(_0574_),
    .B1(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__a31o_1 _1987_ (.A1(\A[8] ),
    .A2(_1061_),
    .A3(_0581_),
    .B1(_0580_),
    .X(_0605_));
 sky130_fd_sc_hd__o211a_1 _1988_ (.A1(\A[11] ),
    .A2(_1064_),
    .B1(_1063_),
    .C1(\A[10] ),
    .X(_0606_));
 sky130_fd_sc_hd__a211o_1 _1989_ (.A1(_0602_),
    .A2(_0605_),
    .B1(_0606_),
    .C1(_0593_),
    .X(_0607_));
 sky130_fd_sc_hd__or3_1 _1990_ (.A(_0601_),
    .B(_0604_),
    .C(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__o21a_1 _1991_ (.A1(_0604_),
    .A2(_0607_),
    .B1(_0601_),
    .X(_0609_));
 sky130_fd_sc_hd__nor2_1 _1992_ (.A(_1149_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__a22o_1 _1993_ (.A1(\A[12] ),
    .A2(_1149_),
    .B1(_0608_),
    .B2(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__o211a_1 _1994_ (.A1(\count[5] ),
    .A2(_0611_),
    .B1(_0422_),
    .C1(_0889_),
    .X(_0211_));
 sky130_fd_sc_hd__xor2_2 _1995_ (.A(\A[13] ),
    .B(_1066_),
    .X(_0612_));
 sky130_fd_sc_hd__o21ai_1 _1996_ (.A1(_0599_),
    .A2(_0609_),
    .B1(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__o311a_1 _1997_ (.A1(_0599_),
    .A2(_0609_),
    .A3(_0612_),
    .B1(_0613_),
    .C1(_1148_),
    .X(_0614_));
 sky130_fd_sc_hd__a21o_1 _1998_ (.A1(\A[13] ),
    .A2(_1149_),
    .B1(\count[5] ),
    .X(_0615_));
 sky130_fd_sc_hd__o221a_1 _1999_ (.A1(\A[12] ),
    .A2(_0873_),
    .B1(_0614_),
    .B2(_0615_),
    .C1(_0889_),
    .X(_0212_));
 sky130_fd_sc_hd__and2_1 _2000_ (.A(\A[14] ),
    .B(_1067_),
    .X(_0616_));
 sky130_fd_sc_hd__nor2_1 _2001_ (.A(\A[14] ),
    .B(_1067_),
    .Y(_0617_));
 sky130_fd_sc_hd__nor2_1 _2002_ (.A(_0616_),
    .B(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__a22o_1 _2003_ (.A1(\A[12] ),
    .A2(_1065_),
    .B1(_1066_),
    .B2(\A[13] ),
    .X(_0619_));
 sky130_fd_sc_hd__o22a_1 _2004_ (.A1(\A[13] ),
    .A2(_1066_),
    .B1(_0609_),
    .B2(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__nand2_1 _2005_ (.A(_0618_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__o21a_1 _2006_ (.A1(_0618_),
    .A2(_0620_),
    .B1(_1148_),
    .X(_0622_));
 sky130_fd_sc_hd__a221o_1 _2007_ (.A1(\A[14] ),
    .A2(_1149_),
    .B1(_0621_),
    .B2(_0622_),
    .C1(\count[5] ),
    .X(_0623_));
 sky130_fd_sc_hd__o211a_1 _2008_ (.A1(\A[13] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0623_),
    .X(_0213_));
 sky130_fd_sc_hd__xor2_1 _2009_ (.A(\A[15] ),
    .B(_1068_),
    .X(_0624_));
 sky130_fd_sc_hd__a21o_1 _2010_ (.A1(_0618_),
    .A2(_0620_),
    .B1(_0616_),
    .X(_0625_));
 sky130_fd_sc_hd__nand2_1 _2011_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__o211a_1 _2012_ (.A1(_0624_),
    .A2(_0625_),
    .B1(_0626_),
    .C1(_1148_),
    .X(_0627_));
 sky130_fd_sc_hd__a21o_1 _2013_ (.A1(\A[15] ),
    .A2(_1149_),
    .B1(\count[5] ),
    .X(_0628_));
 sky130_fd_sc_hd__o221a_1 _2014_ (.A1(\A[14] ),
    .A2(_0873_),
    .B1(_0627_),
    .B2(_0628_),
    .C1(_0889_),
    .X(_0214_));
 sky130_fd_sc_hd__and2_1 _2015_ (.A(_0618_),
    .B(_0624_),
    .X(_0629_));
 sky130_fd_sc_hd__o2111ai_4 _2016_ (.A1(_0604_),
    .A2(_0607_),
    .B1(_0612_),
    .C1(_0629_),
    .D1(_0601_),
    .Y(_0630_));
 sky130_fd_sc_hd__o211a_1 _2017_ (.A1(\A[15] ),
    .A2(_1068_),
    .B1(_1067_),
    .C1(\A[14] ),
    .X(_0631_));
 sky130_fd_sc_hd__o211a_1 _2018_ (.A1(\A[13] ),
    .A2(_1066_),
    .B1(_0619_),
    .C1(_0629_),
    .X(_0632_));
 sky130_fd_sc_hd__a211oi_2 _2019_ (.A1(\A[15] ),
    .A2(_1068_),
    .B1(_0631_),
    .C1(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__and2_1 _2020_ (.A(\A[16] ),
    .B(_1069_),
    .X(_0634_));
 sky130_fd_sc_hd__nor2_1 _2021_ (.A(\A[16] ),
    .B(_1069_),
    .Y(_0635_));
 sky130_fd_sc_hd__or2_1 _2022_ (.A(_0634_),
    .B(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__a21oi_1 _2023_ (.A1(_0630_),
    .A2(_0633_),
    .B1(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__a31o_1 _2024_ (.A1(_0630_),
    .A2(_0633_),
    .A3(_0636_),
    .B1(_1149_),
    .X(_0638_));
 sky130_fd_sc_hd__a2bb2o_1 _2025_ (.A1_N(_0637_),
    .A2_N(_0638_),
    .B1(\A[16] ),
    .B2(_1149_),
    .X(_0639_));
 sky130_fd_sc_hd__o211a_1 _2026_ (.A1(\count[5] ),
    .A2(_0639_),
    .B1(_0442_),
    .C1(_0889_),
    .X(_0215_));
 sky130_fd_sc_hd__and2_1 _2027_ (.A(\A[17] ),
    .B(_1070_),
    .X(_0640_));
 sky130_fd_sc_hd__or2_1 _2028_ (.A(\A[17] ),
    .B(_1070_),
    .X(_0641_));
 sky130_fd_sc_hd__and2b_1 _2029_ (.A_N(_0640_),
    .B(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__or2_1 _2030_ (.A(_0634_),
    .B(_0637_),
    .X(_0643_));
 sky130_fd_sc_hd__xnor2_1 _2031_ (.A(_0642_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__nor2_1 _2032_ (.A(net132),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__a21o_1 _2033_ (.A1(\A[17] ),
    .A2(net132),
    .B1(\count[5] ),
    .X(_0646_));
 sky130_fd_sc_hd__o221a_1 _2034_ (.A1(\A[16] ),
    .A2(_0873_),
    .B1(_0645_),
    .B2(_0646_),
    .C1(_0889_),
    .X(_0216_));
 sky130_fd_sc_hd__and2_1 _2035_ (.A(\A[18] ),
    .B(_1071_),
    .X(_0647_));
 sky130_fd_sc_hd__nor2_1 _2036_ (.A(\A[18] ),
    .B(_1071_),
    .Y(_0648_));
 sky130_fd_sc_hd__nor2_1 _2037_ (.A(_0647_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__a21o_1 _2038_ (.A1(_0641_),
    .A2(_0643_),
    .B1(_0640_),
    .X(_0650_));
 sky130_fd_sc_hd__nand2_1 _2039_ (.A(_0649_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__o21a_1 _2040_ (.A1(_0649_),
    .A2(_0650_),
    .B1(_1148_),
    .X(_0652_));
 sky130_fd_sc_hd__a221o_1 _2041_ (.A1(\A[18] ),
    .A2(net132),
    .B1(_0651_),
    .B2(_0652_),
    .C1(\count[5] ),
    .X(_0653_));
 sky130_fd_sc_hd__o211a_1 _2042_ (.A1(\A[17] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0653_),
    .X(_0217_));
 sky130_fd_sc_hd__xor2_1 _2043_ (.A(\A[19] ),
    .B(_1072_),
    .X(_0654_));
 sky130_fd_sc_hd__a21o_1 _2044_ (.A1(_0649_),
    .A2(_0650_),
    .B1(_0647_),
    .X(_0655_));
 sky130_fd_sc_hd__a21oi_1 _2045_ (.A1(_0654_),
    .A2(_0655_),
    .B1(net132),
    .Y(_0656_));
 sky130_fd_sc_hd__o21a_1 _2046_ (.A1(_0654_),
    .A2(_0655_),
    .B1(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__a21o_1 _2047_ (.A1(\A[19] ),
    .A2(net132),
    .B1(\count[5] ),
    .X(_0658_));
 sky130_fd_sc_hd__o221a_1 _2048_ (.A1(\A[18] ),
    .A2(_0873_),
    .B1(_0657_),
    .B2(_0658_),
    .C1(_0889_),
    .X(_0218_));
 sky130_fd_sc_hd__nand2_1 _2049_ (.A(\A[20] ),
    .B(_1073_),
    .Y(_0659_));
 sky130_fd_sc_hd__or2_1 _2050_ (.A(\A[20] ),
    .B(_1073_),
    .X(_0660_));
 sky130_fd_sc_hd__and2_1 _2051_ (.A(_0659_),
    .B(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__a21o_1 _2052_ (.A1(_0634_),
    .A2(_0641_),
    .B1(_0640_),
    .X(_0662_));
 sky130_fd_sc_hd__and3_1 _2053_ (.A(_0649_),
    .B(_0654_),
    .C(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__o21a_1 _2054_ (.A1(\A[19] ),
    .A2(_1072_),
    .B1(_0647_),
    .X(_0664_));
 sky130_fd_sc_hd__a211oi_2 _2055_ (.A1(\A[19] ),
    .A2(_1072_),
    .B1(_0663_),
    .C1(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand4b_1 _2056_ (.A_N(_0636_),
    .B(_0642_),
    .C(_0649_),
    .D(_0654_),
    .Y(_0666_));
 sky130_fd_sc_hd__a21o_1 _2057_ (.A1(_0630_),
    .A2(_0633_),
    .B1(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__nand2_1 _2058_ (.A(_0665_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__a21bo_1 _2059_ (.A1(_0665_),
    .A2(_0667_),
    .B1_N(_0661_),
    .X(_0669_));
 sky130_fd_sc_hd__o21a_1 _2060_ (.A1(_0661_),
    .A2(_0668_),
    .B1(_1148_),
    .X(_0670_));
 sky130_fd_sc_hd__a221o_1 _2061_ (.A1(\A[20] ),
    .A2(net132),
    .B1(_0669_),
    .B2(_0670_),
    .C1(net134),
    .X(_0671_));
 sky130_fd_sc_hd__o211a_1 _2062_ (.A1(\A[19] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0671_),
    .X(_0219_));
 sky130_fd_sc_hd__and2_1 _2063_ (.A(\A[21] ),
    .B(_1074_),
    .X(_0672_));
 sky130_fd_sc_hd__nor2_1 _2064_ (.A(\A[21] ),
    .B(_1074_),
    .Y(_0673_));
 sky130_fd_sc_hd__nor2_1 _2065_ (.A(_0672_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__and3_1 _2066_ (.A(_0659_),
    .B(_0669_),
    .C(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__a21oi_1 _2067_ (.A1(_0659_),
    .A2(_0669_),
    .B1(_0674_),
    .Y(_0676_));
 sky130_fd_sc_hd__o21a_1 _2068_ (.A1(_0675_),
    .A2(_0676_),
    .B1(_1148_),
    .X(_0677_));
 sky130_fd_sc_hd__a21o_1 _2069_ (.A1(\A[21] ),
    .A2(net132),
    .B1(net134),
    .X(_0678_));
 sky130_fd_sc_hd__o221a_1 _2070_ (.A1(\A[20] ),
    .A2(_0873_),
    .B1(_0677_),
    .B2(_0678_),
    .C1(_0889_),
    .X(_0220_));
 sky130_fd_sc_hd__nand2_1 _2071_ (.A(\A[22] ),
    .B(_1075_),
    .Y(_0679_));
 sky130_fd_sc_hd__or2_1 _2072_ (.A(\A[22] ),
    .B(_1075_),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_1 _2073_ (.A(_0679_),
    .B(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__a21oi_1 _2074_ (.A1(\A[20] ),
    .A2(_1073_),
    .B1(_0672_),
    .Y(_0682_));
 sky130_fd_sc_hd__a21o_1 _2075_ (.A1(_0669_),
    .A2(_0682_),
    .B1(_0673_),
    .X(_0683_));
 sky130_fd_sc_hd__or2_1 _2076_ (.A(_0681_),
    .B(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__a21oi_1 _2077_ (.A1(_0681_),
    .A2(_0683_),
    .B1(net132),
    .Y(_0685_));
 sky130_fd_sc_hd__a221o_1 _2078_ (.A1(\A[22] ),
    .A2(net132),
    .B1(_0684_),
    .B2(_0685_),
    .C1(net134),
    .X(_0686_));
 sky130_fd_sc_hd__o211a_1 _2079_ (.A1(\A[21] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0686_),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_1 _2080_ (.A(\A[23] ),
    .B(_1076_),
    .Y(_0687_));
 sky130_fd_sc_hd__nor2_1 _2081_ (.A(\A[23] ),
    .B(_1076_),
    .Y(_0688_));
 sky130_fd_sc_hd__or2_1 _2082_ (.A(\A[23] ),
    .B(_1076_),
    .X(_0689_));
 sky130_fd_sc_hd__nand2_1 _2083_ (.A(_0687_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__a21oi_1 _2084_ (.A1(_0679_),
    .A2(_0684_),
    .B1(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__a311oi_1 _2085_ (.A1(_0679_),
    .A2(_0684_),
    .A3(_0690_),
    .B1(_0691_),
    .C1(net132),
    .Y(_0692_));
 sky130_fd_sc_hd__a21o_1 _2086_ (.A1(\A[23] ),
    .A2(net132),
    .B1(net134),
    .X(_0693_));
 sky130_fd_sc_hd__o221a_1 _2087_ (.A1(\A[22] ),
    .A2(_0873_),
    .B1(_0692_),
    .B2(_0693_),
    .C1(_0889_),
    .X(_0222_));
 sky130_fd_sc_hd__nand2_1 _2088_ (.A(\A[24] ),
    .B(_1077_),
    .Y(_0694_));
 sky130_fd_sc_hd__or2_1 _2089_ (.A(\A[24] ),
    .B(_1077_),
    .X(_0695_));
 sky130_fd_sc_hd__nand2_1 _2090_ (.A(_0694_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__or2_1 _2091_ (.A(_0681_),
    .B(_0690_),
    .X(_0697_));
 sky130_fd_sc_hd__nand2_1 _2092_ (.A(_0661_),
    .B(_0674_),
    .Y(_0698_));
 sky130_fd_sc_hd__o22a_1 _2093_ (.A1(_0673_),
    .A2(_0682_),
    .B1(_0698_),
    .B2(_0665_),
    .X(_0699_));
 sky130_fd_sc_hd__o221a_1 _2094_ (.A1(_0679_),
    .A2(_0688_),
    .B1(_0697_),
    .B2(_0699_),
    .C1(_0687_),
    .X(_0700_));
 sky130_fd_sc_hd__a2111o_1 _2095_ (.A1(_0630_),
    .A2(_0633_),
    .B1(_0666_),
    .C1(_0697_),
    .D1(_0698_),
    .X(_0701_));
 sky130_fd_sc_hd__a21o_1 _2096_ (.A1(_0700_),
    .A2(_0701_),
    .B1(_0696_),
    .X(_0702_));
 sky130_fd_sc_hd__a31oi_1 _2097_ (.A1(_0696_),
    .A2(_0700_),
    .A3(_0701_),
    .B1(net132),
    .Y(_0703_));
 sky130_fd_sc_hd__a221o_1 _2098_ (.A1(\A[24] ),
    .A2(net132),
    .B1(_0702_),
    .B2(_0703_),
    .C1(net134),
    .X(_0704_));
 sky130_fd_sc_hd__o211a_1 _2099_ (.A1(\A[23] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0704_),
    .X(_0223_));
 sky130_fd_sc_hd__nor2_1 _2100_ (.A(\A[25] ),
    .B(_1078_),
    .Y(_0705_));
 sky130_fd_sc_hd__and2_1 _2101_ (.A(\A[25] ),
    .B(_1078_),
    .X(_0706_));
 sky130_fd_sc_hd__or2_1 _2102_ (.A(_0705_),
    .B(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__a21oi_1 _2103_ (.A1(_0694_),
    .A2(_0702_),
    .B1(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__a311oi_1 _2104_ (.A1(_0694_),
    .A2(_0702_),
    .A3(_0707_),
    .B1(_0708_),
    .C1(net132),
    .Y(_0709_));
 sky130_fd_sc_hd__a21o_1 _2105_ (.A1(\A[25] ),
    .A2(net132),
    .B1(net134),
    .X(_0710_));
 sky130_fd_sc_hd__o211a_1 _2106_ (.A1(_0709_),
    .A2(_0710_),
    .B1(_0889_),
    .C1(_0483_),
    .X(_0224_));
 sky130_fd_sc_hd__nand2_1 _2107_ (.A(\A[26] ),
    .B(_1079_),
    .Y(_0711_));
 sky130_fd_sc_hd__or2_1 _2108_ (.A(\A[26] ),
    .B(_1079_),
    .X(_0712_));
 sky130_fd_sc_hd__nand2_1 _2109_ (.A(_0711_),
    .B(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__a21oi_1 _2110_ (.A1(\A[24] ),
    .A2(_1077_),
    .B1(_0706_),
    .Y(_0714_));
 sky130_fd_sc_hd__a21o_1 _2111_ (.A1(_0702_),
    .A2(_0714_),
    .B1(_0705_),
    .X(_0715_));
 sky130_fd_sc_hd__or2_1 _2112_ (.A(_0713_),
    .B(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__a21oi_1 _2113_ (.A1(_0713_),
    .A2(_0715_),
    .B1(net132),
    .Y(_0717_));
 sky130_fd_sc_hd__a221o_1 _2114_ (.A1(\A[26] ),
    .A2(net132),
    .B1(_0716_),
    .B2(_0717_),
    .C1(net134),
    .X(_0718_));
 sky130_fd_sc_hd__o211a_1 _2115_ (.A1(\A[25] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0718_),
    .X(_0225_));
 sky130_fd_sc_hd__nand2_1 _2116_ (.A(\A[27] ),
    .B(_1080_),
    .Y(_0719_));
 sky130_fd_sc_hd__or2_1 _2117_ (.A(\A[27] ),
    .B(_1080_),
    .X(_0720_));
 sky130_fd_sc_hd__nand2_1 _2118_ (.A(_0719_),
    .B(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__a21oi_1 _2119_ (.A1(_0711_),
    .A2(_0716_),
    .B1(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__a311oi_1 _2120_ (.A1(_0711_),
    .A2(_0716_),
    .A3(_0721_),
    .B1(_0722_),
    .C1(net132),
    .Y(_0723_));
 sky130_fd_sc_hd__a21o_1 _2121_ (.A1(\A[27] ),
    .A2(net132),
    .B1(net134),
    .X(_0724_));
 sky130_fd_sc_hd__o221a_1 _2122_ (.A1(\A[26] ),
    .A2(_0873_),
    .B1(_0723_),
    .B2(_0724_),
    .C1(_0889_),
    .X(_0226_));
 sky130_fd_sc_hd__or2_1 _2123_ (.A(_0713_),
    .B(_0721_),
    .X(_0725_));
 sky130_fd_sc_hd__or3_1 _2124_ (.A(_0696_),
    .B(_0707_),
    .C(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__a21o_1 _2125_ (.A1(_0700_),
    .A2(_0701_),
    .B1(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__o21bai_1 _2126_ (.A1(\A[27] ),
    .A2(_1080_),
    .B1_N(_0711_),
    .Y(_0728_));
 sky130_fd_sc_hd__o311a_1 _2127_ (.A1(_0705_),
    .A2(_0714_),
    .A3(_0725_),
    .B1(_0728_),
    .C1(_0719_),
    .X(_0729_));
 sky130_fd_sc_hd__nand2_1 _2128_ (.A(\A[28] ),
    .B(_1081_),
    .Y(_0730_));
 sky130_fd_sc_hd__or2_1 _2129_ (.A(\A[28] ),
    .B(_1081_),
    .X(_0731_));
 sky130_fd_sc_hd__nand2_1 _2130_ (.A(_0730_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__a21o_1 _2131_ (.A1(_0727_),
    .A2(_0729_),
    .B1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__a31oi_1 _2132_ (.A1(_0727_),
    .A2(_0729_),
    .A3(_0732_),
    .B1(net132),
    .Y(_0734_));
 sky130_fd_sc_hd__a221o_1 _2133_ (.A1(\A[28] ),
    .A2(net132),
    .B1(_0733_),
    .B2(_0734_),
    .C1(net134),
    .X(_0735_));
 sky130_fd_sc_hd__o211a_1 _2134_ (.A1(\A[27] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0735_),
    .X(_0227_));
 sky130_fd_sc_hd__nand2_1 _2135_ (.A(\A[29] ),
    .B(_1082_),
    .Y(_0736_));
 sky130_fd_sc_hd__or2_1 _2136_ (.A(\A[29] ),
    .B(_1082_),
    .X(_0737_));
 sky130_fd_sc_hd__inv_2 _2137_ (.A(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__nand2_1 _2138_ (.A(_0736_),
    .B(_0737_),
    .Y(_0739_));
 sky130_fd_sc_hd__nand2_1 _2139_ (.A(_0730_),
    .B(_0733_),
    .Y(_0740_));
 sky130_fd_sc_hd__a31o_1 _2140_ (.A1(_0730_),
    .A2(_0733_),
    .A3(_0739_),
    .B1(net132),
    .X(_0741_));
 sky130_fd_sc_hd__a31oi_1 _2141_ (.A1(_0736_),
    .A2(_0737_),
    .A3(_0740_),
    .B1(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__a21o_1 _2142_ (.A1(\A[29] ),
    .A2(net132),
    .B1(net134),
    .X(_0743_));
 sky130_fd_sc_hd__o221a_1 _2143_ (.A1(\A[28] ),
    .A2(_0873_),
    .B1(_0742_),
    .B2(_0743_),
    .C1(_0889_),
    .X(_0228_));
 sky130_fd_sc_hd__or2_1 _2144_ (.A(\A[30] ),
    .B(_1083_),
    .X(_0744_));
 sky130_fd_sc_hd__and2_1 _2145_ (.A(\A[30] ),
    .B(_1083_),
    .X(_0745_));
 sky130_fd_sc_hd__nand2_1 _2146_ (.A(\A[30] ),
    .B(_1083_),
    .Y(_0746_));
 sky130_fd_sc_hd__nand2_1 _2147_ (.A(_0744_),
    .B(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__nand2_1 _2148_ (.A(_0730_),
    .B(_0736_),
    .Y(_0748_));
 sky130_fd_sc_hd__inv_2 _2149_ (.A(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__nand2_1 _2150_ (.A(_0737_),
    .B(_0740_),
    .Y(_0750_));
 sky130_fd_sc_hd__a211oi_1 _2151_ (.A1(_0733_),
    .A2(_0749_),
    .B1(_0747_),
    .C1(_0738_),
    .Y(_0751_));
 sky130_fd_sc_hd__a311oi_1 _2152_ (.A1(_0736_),
    .A2(_0747_),
    .A3(_0750_),
    .B1(_0751_),
    .C1(net132),
    .Y(_0752_));
 sky130_fd_sc_hd__a21o_1 _2153_ (.A1(\A[30] ),
    .A2(net132),
    .B1(net134),
    .X(_0753_));
 sky130_fd_sc_hd__o221a_1 _2154_ (.A1(\A[29] ),
    .A2(_0873_),
    .B1(_0752_),
    .B2(_0753_),
    .C1(_0889_),
    .X(_0229_));
 sky130_fd_sc_hd__or2_1 _2155_ (.A(\A[31] ),
    .B(_1084_),
    .X(_0754_));
 sky130_fd_sc_hd__nand2_1 _2156_ (.A(\A[31] ),
    .B(_1084_),
    .Y(_0755_));
 sky130_fd_sc_hd__nand2_1 _2157_ (.A(_0754_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__inv_2 _2158_ (.A(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__o21ai_1 _2159_ (.A1(_0745_),
    .A2(_0751_),
    .B1(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__o31a_1 _2160_ (.A1(_0745_),
    .A2(_0751_),
    .A3(_0757_),
    .B1(_1148_),
    .X(_0759_));
 sky130_fd_sc_hd__a221o_1 _2161_ (.A1(\A[31] ),
    .A2(net132),
    .B1(_0758_),
    .B2(_0759_),
    .C1(net134),
    .X(_0760_));
 sky130_fd_sc_hd__o211a_1 _2162_ (.A1(\A[30] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0760_),
    .X(_0230_));
 sky130_fd_sc_hd__or4_1 _2163_ (.A(_0732_),
    .B(_0739_),
    .C(_0747_),
    .D(_0756_),
    .X(_0761_));
 sky130_fd_sc_hd__a21oi_2 _2164_ (.A1(_0727_),
    .A2(_0729_),
    .B1(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__a21o_1 _2165_ (.A1(_0727_),
    .A2(_0729_),
    .B1(_0761_),
    .X(_0763_));
 sky130_fd_sc_hd__a21bo_1 _2166_ (.A1(_0746_),
    .A2(_0755_),
    .B1_N(_0754_),
    .X(_0764_));
 sky130_fd_sc_hd__o41a_2 _2167_ (.A1(_0738_),
    .A2(_0747_),
    .A3(_0749_),
    .A4(_0756_),
    .B1(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__inv_2 _2168_ (.A(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__a21oi_2 _2169_ (.A1(_0763_),
    .A2(_0765_),
    .B1(net132),
    .Y(_0767_));
 sky130_fd_sc_hd__nand2_1 _2170_ (.A(\A[32] ),
    .B(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__or2_1 _2171_ (.A(\A[32] ),
    .B(_0767_),
    .X(_0769_));
 sky130_fd_sc_hd__a21o_1 _2172_ (.A1(_0768_),
    .A2(_0769_),
    .B1(net135),
    .X(_0770_));
 sky130_fd_sc_hd__o211a_1 _2173_ (.A1(\A[31] ),
    .A2(_0873_),
    .B1(_0889_),
    .C1(_0770_),
    .X(_0231_));
 sky130_fd_sc_hd__a31o_1 _2174_ (.A1(\A[33] ),
    .A2(\A[32] ),
    .A3(_0767_),
    .B1(net135),
    .X(_0771_));
 sky130_fd_sc_hd__a21oi_1 _2175_ (.A1(\A[32] ),
    .A2(_0767_),
    .B1(\A[33] ),
    .Y(_0772_));
 sky130_fd_sc_hd__o2bb2a_1 _2176_ (.A1_N(\A[32] ),
    .A2_N(net135),
    .B1(_0771_),
    .B2(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__nor2_1 _2177_ (.A(net66),
    .B(_0773_),
    .Y(_0232_));
 sky130_fd_sc_hd__nand2_1 _2178_ (.A(\A[33] ),
    .B(net135),
    .Y(_0774_));
 sky130_fd_sc_hd__a41o_1 _2179_ (.A1(\A[33] ),
    .A2(\A[32] ),
    .A3(_0873_),
    .A4(_0767_),
    .B1(\A[34] ),
    .X(_0775_));
 sky130_fd_sc_hd__a21bo_1 _2180_ (.A1(\A[34] ),
    .A2(_0771_),
    .B1_N(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__a21oi_1 _2181_ (.A1(_0774_),
    .A2(_0776_),
    .B1(net66),
    .Y(_0233_));
 sky130_fd_sc_hd__a22o_1 _2182_ (.A1(\A[35] ),
    .A2(_0873_),
    .B1(_0771_),
    .B2(\A[34] ),
    .X(_0777_));
 sky130_fd_sc_hd__and4_1 _2183_ (.A(\A[35] ),
    .B(\A[34] ),
    .C(\A[33] ),
    .D(\A[32] ),
    .X(_0778_));
 sky130_fd_sc_hd__o2111ai_2 _2184_ (.A1(_0762_),
    .A2(_0766_),
    .B1(_0778_),
    .C1(_1148_),
    .D1(_0873_),
    .Y(_0779_));
 sky130_fd_sc_hd__and3_1 _2185_ (.A(_0889_),
    .B(_0777_),
    .C(_0779_),
    .X(_0234_));
 sky130_fd_sc_hd__nand2_1 _2186_ (.A(\A[35] ),
    .B(net135),
    .Y(_0780_));
 sky130_fd_sc_hd__a21o_1 _2187_ (.A1(_0767_),
    .A2(_0778_),
    .B1(net135),
    .X(_0781_));
 sky130_fd_sc_hd__mux2_1 _2188_ (.A0(_0779_),
    .A1(_0781_),
    .S(\A[36] ),
    .X(_0782_));
 sky130_fd_sc_hd__a21oi_1 _2189_ (.A1(_0780_),
    .A2(_0782_),
    .B1(net66),
    .Y(_0235_));
 sky130_fd_sc_hd__a22oi_1 _2190_ (.A1(\A[37] ),
    .A2(_0873_),
    .B1(_0781_),
    .B2(\A[36] ),
    .Y(_0783_));
 sky130_fd_sc_hd__and2_1 _2191_ (.A(\A[37] ),
    .B(\A[36] ),
    .X(_0784_));
 sky130_fd_sc_hd__and2b_1 _2192_ (.A_N(_0779_),
    .B(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__nor3_1 _2193_ (.A(net66),
    .B(_0783_),
    .C(_0785_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _2194_ (.A(\A[37] ),
    .B(net135),
    .Y(_0786_));
 sky130_fd_sc_hd__o21a_1 _2195_ (.A1(net135),
    .A2(_0784_),
    .B1(\A[38] ),
    .X(_0787_));
 sky130_fd_sc_hd__a2bb2o_1 _2196_ (.A1_N(\A[38] ),
    .A2_N(_0785_),
    .B1(_0787_),
    .B2(_0781_),
    .X(_0788_));
 sky130_fd_sc_hd__a21oi_1 _2197_ (.A1(_0786_),
    .A2(_0788_),
    .B1(net66),
    .Y(_0237_));
 sky130_fd_sc_hd__a22o_1 _2198_ (.A1(\A[39] ),
    .A2(_0873_),
    .B1(_0781_),
    .B2(_0787_),
    .X(_0789_));
 sky130_fd_sc_hd__and3_1 _2199_ (.A(\A[39] ),
    .B(\A[38] ),
    .C(_0784_),
    .X(_0790_));
 sky130_fd_sc_hd__nand2b_1 _2200_ (.A_N(_0779_),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__and4_1 _2201_ (.A(\A[39] ),
    .B(\A[38] ),
    .C(_0778_),
    .D(_0784_),
    .X(_0792_));
 sky130_fd_sc_hd__and3_1 _2202_ (.A(_0889_),
    .B(_0789_),
    .C(_0791_),
    .X(_0238_));
 sky130_fd_sc_hd__nand2_1 _2203_ (.A(\A[39] ),
    .B(net135),
    .Y(_0793_));
 sky130_fd_sc_hd__o2111a_1 _2204_ (.A1(_0762_),
    .A2(_0766_),
    .B1(_0778_),
    .C1(_0790_),
    .D1(_1148_),
    .X(_0794_));
 sky130_fd_sc_hd__or2_1 _2205_ (.A(net135),
    .B(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _2206_ (.A0(_0791_),
    .A1(_0795_),
    .S(\A[40] ),
    .X(_0796_));
 sky130_fd_sc_hd__a21oi_1 _2207_ (.A1(_0793_),
    .A2(_0796_),
    .B1(net66),
    .Y(_0239_));
 sky130_fd_sc_hd__a22o_1 _2208_ (.A1(\A[41] ),
    .A2(_0873_),
    .B1(_0795_),
    .B2(\A[40] ),
    .X(_0797_));
 sky130_fd_sc_hd__and2_1 _2209_ (.A(\A[41] ),
    .B(\A[40] ),
    .X(_0798_));
 sky130_fd_sc_hd__nand2_1 _2210_ (.A(\A[41] ),
    .B(\A[40] ),
    .Y(_0799_));
 sky130_fd_sc_hd__o211a_1 _2211_ (.A1(_0791_),
    .A2(_0799_),
    .B1(_0797_),
    .C1(_0889_),
    .X(_0240_));
 sky130_fd_sc_hd__nand2_1 _2212_ (.A(\A[41] ),
    .B(net135),
    .Y(_0800_));
 sky130_fd_sc_hd__a21o_1 _2213_ (.A1(_0794_),
    .A2(_0798_),
    .B1(net135),
    .X(_0801_));
 sky130_fd_sc_hd__a31o_1 _2214_ (.A1(_0873_),
    .A2(_0794_),
    .A3(_0798_),
    .B1(\A[42] ),
    .X(_0802_));
 sky130_fd_sc_hd__a21bo_1 _2215_ (.A1(\A[42] ),
    .A2(_0801_),
    .B1_N(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__a21oi_1 _2216_ (.A1(_0800_),
    .A2(_0803_),
    .B1(net66),
    .Y(_0241_));
 sky130_fd_sc_hd__a22o_1 _2217_ (.A1(\A[43] ),
    .A2(_0873_),
    .B1(_0801_),
    .B2(\A[42] ),
    .X(_0804_));
 sky130_fd_sc_hd__and3_1 _2218_ (.A(\A[43] ),
    .B(\A[42] ),
    .C(_0798_),
    .X(_0805_));
 sky130_fd_sc_hd__o2111a_1 _2219_ (.A1(_0762_),
    .A2(_0766_),
    .B1(_0792_),
    .C1(_0805_),
    .D1(_1148_),
    .X(_0806_));
 sky130_fd_sc_hd__nand2_1 _2220_ (.A(_0873_),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__and3_1 _2221_ (.A(_0889_),
    .B(_0804_),
    .C(_0807_),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_1 _2222_ (.A(\A[43] ),
    .B(net135),
    .Y(_0808_));
 sky130_fd_sc_hd__or2_1 _2223_ (.A(net135),
    .B(_0806_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _2224_ (.A0(_0807_),
    .A1(_0809_),
    .S(\A[44] ),
    .X(_0810_));
 sky130_fd_sc_hd__a21oi_1 _2225_ (.A1(_0808_),
    .A2(_0810_),
    .B1(net66),
    .Y(_0243_));
 sky130_fd_sc_hd__a22oi_1 _2226_ (.A1(\A[45] ),
    .A2(_0873_),
    .B1(_0809_),
    .B2(\A[44] ),
    .Y(_0811_));
 sky130_fd_sc_hd__and2_1 _2227_ (.A(\A[45] ),
    .B(\A[44] ),
    .X(_0812_));
 sky130_fd_sc_hd__and3_1 _2228_ (.A(_0873_),
    .B(_0806_),
    .C(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__nor3_1 _2229_ (.A(net66),
    .B(_0811_),
    .C(_0813_),
    .Y(_0244_));
 sky130_fd_sc_hd__nand2_1 _2230_ (.A(\A[45] ),
    .B(net135),
    .Y(_0814_));
 sky130_fd_sc_hd__o21a_1 _2231_ (.A1(net135),
    .A2(_0812_),
    .B1(\A[46] ),
    .X(_0815_));
 sky130_fd_sc_hd__a2bb2o_1 _2232_ (.A1_N(\A[46] ),
    .A2_N(_0813_),
    .B1(_0815_),
    .B2(_0809_),
    .X(_0816_));
 sky130_fd_sc_hd__a21oi_1 _2233_ (.A1(_0814_),
    .A2(_0816_),
    .B1(net66),
    .Y(_0245_));
 sky130_fd_sc_hd__a22o_1 _2234_ (.A1(\A[47] ),
    .A2(_0873_),
    .B1(_0809_),
    .B2(_0815_),
    .X(_0817_));
 sky130_fd_sc_hd__and3_1 _2235_ (.A(\A[47] ),
    .B(\A[46] ),
    .C(_0812_),
    .X(_0818_));
 sky130_fd_sc_hd__and4_1 _2236_ (.A(_0778_),
    .B(_0790_),
    .C(_0805_),
    .D(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__inv_2 _2237_ (.A(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__a2111o_2 _2238_ (.A1(_0763_),
    .A2(_0765_),
    .B1(_0820_),
    .C1(net132),
    .D1(net134),
    .X(_0821_));
 sky130_fd_sc_hd__and3_1 _2239_ (.A(_0792_),
    .B(_0805_),
    .C(_0818_),
    .X(_0822_));
 sky130_fd_sc_hd__and3_1 _2240_ (.A(_0889_),
    .B(_0817_),
    .C(_0821_),
    .X(_0246_));
 sky130_fd_sc_hd__nand2_1 _2241_ (.A(\A[47] ),
    .B(net135),
    .Y(_0823_));
 sky130_fd_sc_hd__a21o_2 _2242_ (.A1(_0767_),
    .A2(_0822_),
    .B1(net134),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _2243_ (.A0(_0821_),
    .A1(_0824_),
    .S(\A[48] ),
    .X(_0825_));
 sky130_fd_sc_hd__a21oi_1 _2244_ (.A1(_0823_),
    .A2(_0825_),
    .B1(net66),
    .Y(_0247_));
 sky130_fd_sc_hd__a22oi_1 _2245_ (.A1(\A[49] ),
    .A2(_0873_),
    .B1(_0824_),
    .B2(\A[48] ),
    .Y(_0826_));
 sky130_fd_sc_hd__and2_1 _2246_ (.A(\A[49] ),
    .B(\A[48] ),
    .X(_0827_));
 sky130_fd_sc_hd__and2b_1 _2247_ (.A_N(_0821_),
    .B(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__nor3_1 _2248_ (.A(net66),
    .B(_0826_),
    .C(_0828_),
    .Y(_0248_));
 sky130_fd_sc_hd__nand2_1 _2249_ (.A(\A[49] ),
    .B(net134),
    .Y(_0829_));
 sky130_fd_sc_hd__o21a_1 _2250_ (.A1(net134),
    .A2(_0827_),
    .B1(\A[50] ),
    .X(_0830_));
 sky130_fd_sc_hd__a2bb2o_1 _2251_ (.A1_N(\A[50] ),
    .A2_N(_0828_),
    .B1(_0830_),
    .B2(_0824_),
    .X(_0831_));
 sky130_fd_sc_hd__a21oi_1 _2252_ (.A1(_0829_),
    .A2(_0831_),
    .B1(net66),
    .Y(_0249_));
 sky130_fd_sc_hd__a22o_1 _2253_ (.A1(\A[51] ),
    .A2(_0873_),
    .B1(_0824_),
    .B2(_0830_),
    .X(_0832_));
 sky130_fd_sc_hd__and3_1 _2254_ (.A(\A[51] ),
    .B(\A[50] ),
    .C(_0827_),
    .X(_0833_));
 sky130_fd_sc_hd__nand3_1 _2255_ (.A(\A[51] ),
    .B(\A[50] ),
    .C(_0827_),
    .Y(_0834_));
 sky130_fd_sc_hd__o211a_1 _2256_ (.A1(_0821_),
    .A2(_0834_),
    .B1(_0832_),
    .C1(_0889_),
    .X(_0250_));
 sky130_fd_sc_hd__nand2_1 _2257_ (.A(\A[51] ),
    .B(\count[5] ),
    .Y(_0835_));
 sky130_fd_sc_hd__nand2_1 _2258_ (.A(_0873_),
    .B(_0834_),
    .Y(_0836_));
 sky130_fd_sc_hd__o21ba_1 _2259_ (.A1(_0821_),
    .A2(_0834_),
    .B1_N(\A[52] ),
    .X(_0837_));
 sky130_fd_sc_hd__a31o_1 _2260_ (.A1(\A[52] ),
    .A2(_0824_),
    .A3(_0836_),
    .B1(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__a21oi_1 _2261_ (.A1(_0835_),
    .A2(_0838_),
    .B1(net66),
    .Y(_0251_));
 sky130_fd_sc_hd__a32o_1 _2262_ (.A1(\A[52] ),
    .A2(_0824_),
    .A3(_0836_),
    .B1(_0873_),
    .B2(\A[53] ),
    .X(_0839_));
 sky130_fd_sc_hd__and2_1 _2263_ (.A(\A[53] ),
    .B(\A[52] ),
    .X(_0840_));
 sky130_fd_sc_hd__or3b_1 _2264_ (.A(_0821_),
    .B(_0834_),
    .C_N(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__and3_1 _2265_ (.A(_0889_),
    .B(_0839_),
    .C(_0841_),
    .X(_0252_));
 sky130_fd_sc_hd__nand2_1 _2266_ (.A(\A[53] ),
    .B(net135),
    .Y(_0842_));
 sky130_fd_sc_hd__o21a_1 _2267_ (.A1(net134),
    .A2(_0840_),
    .B1(\A[54] ),
    .X(_0843_));
 sky130_fd_sc_hd__a32o_1 _2268_ (.A1(_0824_),
    .A2(_0836_),
    .A3(_0843_),
    .B1(_0841_),
    .B2(_0871_),
    .X(_0844_));
 sky130_fd_sc_hd__a21oi_1 _2269_ (.A1(_0842_),
    .A2(_0844_),
    .B1(net66),
    .Y(_0253_));
 sky130_fd_sc_hd__a32o_1 _2270_ (.A1(_0824_),
    .A2(_0836_),
    .A3(_0843_),
    .B1(_0873_),
    .B2(\A[55] ),
    .X(_0845_));
 sky130_fd_sc_hd__and4_1 _2271_ (.A(\A[55] ),
    .B(\A[54] ),
    .C(_0833_),
    .D(_0840_),
    .X(_0846_));
 sky130_fd_sc_hd__nand4_1 _2272_ (.A(\A[55] ),
    .B(\A[54] ),
    .C(_0833_),
    .D(_0840_),
    .Y(_0847_));
 sky130_fd_sc_hd__o2111a_1 _2273_ (.A1(_0762_),
    .A2(_0766_),
    .B1(_0822_),
    .C1(_0846_),
    .D1(_1148_),
    .X(_0848_));
 sky130_fd_sc_hd__o211a_1 _2274_ (.A1(_0821_),
    .A2(_0847_),
    .B1(_0845_),
    .C1(_0889_),
    .X(_0254_));
 sky130_fd_sc_hd__a2111o_1 _2275_ (.A1(_0763_),
    .A2(_0765_),
    .B1(_0820_),
    .C1(_0847_),
    .D1(_1149_),
    .X(_0849_));
 sky130_fd_sc_hd__o21a_1 _2276_ (.A1(net135),
    .A2(_0848_),
    .B1(\A[56] ),
    .X(_0850_));
 sky130_fd_sc_hd__a21oi_1 _2277_ (.A1(_0873_),
    .A2(_0848_),
    .B1(\A[56] ),
    .Y(_0851_));
 sky130_fd_sc_hd__o2bb2a_1 _2278_ (.A1_N(\A[55] ),
    .A2_N(net135),
    .B1(_0850_),
    .B2(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__nor2_1 _2279_ (.A(net66),
    .B(_0852_),
    .Y(_0255_));
 sky130_fd_sc_hd__a21o_1 _2280_ (.A1(\A[57] ),
    .A2(_0873_),
    .B1(_0850_),
    .X(_0853_));
 sky130_fd_sc_hd__nand2_1 _2281_ (.A(\A[57] ),
    .B(\A[56] ),
    .Y(_0854_));
 sky130_fd_sc_hd__or3_1 _2282_ (.A(net135),
    .B(_0849_),
    .C(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__and3_1 _2283_ (.A(_0889_),
    .B(_0853_),
    .C(_0855_),
    .X(_0256_));
 sky130_fd_sc_hd__nand2_1 _2284_ (.A(\A[57] ),
    .B(net135),
    .Y(_0856_));
 sky130_fd_sc_hd__o21ai_1 _2285_ (.A1(_0849_),
    .A2(_0854_),
    .B1(_0873_),
    .Y(_0857_));
 sky130_fd_sc_hd__mux2_1 _2286_ (.A0(_0855_),
    .A1(_0857_),
    .S(\A[58] ),
    .X(_0858_));
 sky130_fd_sc_hd__a21oi_1 _2287_ (.A1(_0856_),
    .A2(_0858_),
    .B1(net66),
    .Y(_0257_));
 sky130_fd_sc_hd__a22o_1 _2288_ (.A1(\A[59] ),
    .A2(_0873_),
    .B1(_0857_),
    .B2(\A[58] ),
    .X(_0859_));
 sky130_fd_sc_hd__nand2_1 _2289_ (.A(\A[59] ),
    .B(\A[58] ),
    .Y(_0860_));
 sky130_fd_sc_hd__nor2_1 _2290_ (.A(_0854_),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__or4_1 _2291_ (.A(net135),
    .B(_0849_),
    .C(_0854_),
    .D(_0860_),
    .X(_0862_));
 sky130_fd_sc_hd__and3_1 _2292_ (.A(_0889_),
    .B(_0859_),
    .C(_0862_),
    .X(_0258_));
 sky130_fd_sc_hd__nand2_1 _2293_ (.A(\A[59] ),
    .B(net135),
    .Y(_0863_));
 sky130_fd_sc_hd__a21o_1 _2294_ (.A1(_0848_),
    .A2(_0861_),
    .B1(net135),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _2295_ (.A0(_0862_),
    .A1(_0864_),
    .S(\A[60] ),
    .X(_0865_));
 sky130_fd_sc_hd__a21oi_1 _2296_ (.A1(_0863_),
    .A2(_0865_),
    .B1(net66),
    .Y(_0259_));
 sky130_fd_sc_hd__o2bb2a_1 _2297_ (.A1_N(_0864_),
    .A2_N(\A[60] ),
    .B1(_0870_),
    .B2(net135),
    .X(_0866_));
 sky130_fd_sc_hd__and4_1 _2298_ (.A(\A[61] ),
    .B(\A[60] ),
    .C(_0848_),
    .D(_0861_),
    .X(_0867_));
 sky130_fd_sc_hd__a211oi_1 _2299_ (.A1(_0873_),
    .A2(_0867_),
    .B1(_0866_),
    .C1(net66),
    .Y(_0260_));
 sky130_fd_sc_hd__nand2_1 _2300_ (.A(_0870_),
    .B(net135),
    .Y(_0868_));
 sky130_fd_sc_hd__xor2_1 _2301_ (.A(\A[62] ),
    .B(_0867_),
    .X(_0869_));
 sky130_fd_sc_hd__o211a_1 _2302_ (.A1(net135),
    .A2(_0869_),
    .B1(_0868_),
    .C1(_0889_),
    .X(_0261_));
 sky130_fd_sc_hd__o211a_1 _2303_ (.A1(net135),
    .A2(_0867_),
    .B1(_0889_),
    .C1(\A[62] ),
    .X(_0262_));
 sky130_fd_sc_hd__dfxtp_4 _2304_ (.CLK(net1),
    .D(_0000_),
    .Q(sign));
 sky130_fd_sc_hd__dfxtp_1 _2305_ (.CLK(net1),
    .D(_0001_),
    .Q(\abs_multiplier[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2306_ (.CLK(net1),
    .D(_0002_),
    .Q(\abs_multiplier[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2307_ (.CLK(net1),
    .D(_0003_),
    .Q(\abs_multiplier[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2308_ (.CLK(net1),
    .D(_0004_),
    .Q(\abs_multiplier[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2309_ (.CLK(net1),
    .D(_0005_),
    .Q(\abs_multiplier[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2310_ (.CLK(net1),
    .D(_0006_),
    .Q(\abs_multiplier[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2311_ (.CLK(net1),
    .D(_0007_),
    .Q(\abs_multiplier[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2312_ (.CLK(net1),
    .D(_0008_),
    .Q(\abs_multiplier[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2313_ (.CLK(net1),
    .D(_0009_),
    .Q(\abs_multiplier[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2314_ (.CLK(net1),
    .D(_0010_),
    .Q(\abs_multiplier[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2315_ (.CLK(net1),
    .D(_0011_),
    .Q(\abs_multiplier[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2316_ (.CLK(net1),
    .D(_0012_),
    .Q(\abs_multiplier[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2317_ (.CLK(net1),
    .D(_0013_),
    .Q(\abs_multiplier[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2318_ (.CLK(net1),
    .D(_0014_),
    .Q(\abs_multiplier[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2319_ (.CLK(net1),
    .D(_0015_),
    .Q(\abs_multiplier[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2320_ (.CLK(net1),
    .D(_0016_),
    .Q(\abs_multiplier[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2321_ (.CLK(net1),
    .D(_0017_),
    .Q(\abs_multiplier[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2322_ (.CLK(net1),
    .D(_0018_),
    .Q(\abs_multiplier[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2323_ (.CLK(net1),
    .D(_0019_),
    .Q(\abs_multiplier[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2324_ (.CLK(net1),
    .D(_0020_),
    .Q(\abs_multiplier[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2325_ (.CLK(net1),
    .D(_0021_),
    .Q(\abs_multiplier[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2326_ (.CLK(net1),
    .D(_0022_),
    .Q(\abs_multiplier[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2327_ (.CLK(net1),
    .D(_0023_),
    .Q(\abs_multiplier[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2328_ (.CLK(net1),
    .D(_0024_),
    .Q(\abs_multiplier[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2329_ (.CLK(net1),
    .D(_0025_),
    .Q(\abs_multiplier[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2330_ (.CLK(net1),
    .D(_0026_),
    .Q(\abs_multiplier[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2331_ (.CLK(net1),
    .D(_0027_),
    .Q(\abs_multiplier[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2332_ (.CLK(net1),
    .D(_0028_),
    .Q(\abs_multiplier[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2333_ (.CLK(net1),
    .D(_0029_),
    .Q(\abs_multiplier[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2334_ (.CLK(net1),
    .D(_0030_),
    .Q(\abs_multiplier[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2335_ (.CLK(net1),
    .D(_0031_),
    .Q(\abs_multiplier[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2336_ (.CLK(net1),
    .D(_0032_),
    .Q(\abs_multiplicand[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2337_ (.CLK(net1),
    .D(_0033_),
    .Q(\abs_multiplicand[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2338_ (.CLK(net1),
    .D(_0034_),
    .Q(\abs_multiplicand[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2339_ (.CLK(net1),
    .D(_0035_),
    .Q(\abs_multiplicand[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2340_ (.CLK(net1),
    .D(_0036_),
    .Q(\abs_multiplicand[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2341_ (.CLK(net1),
    .D(_0037_),
    .Q(\abs_multiplicand[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2342_ (.CLK(net1),
    .D(_0038_),
    .Q(\abs_multiplicand[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2343_ (.CLK(net1),
    .D(_0039_),
    .Q(\abs_multiplicand[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2344_ (.CLK(net1),
    .D(_0040_),
    .Q(\abs_multiplicand[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2345_ (.CLK(net1),
    .D(_0041_),
    .Q(\abs_multiplicand[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2346_ (.CLK(net1),
    .D(_0042_),
    .Q(\abs_multiplicand[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2347_ (.CLK(net1),
    .D(_0043_),
    .Q(\abs_multiplicand[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2348_ (.CLK(net1),
    .D(_0044_),
    .Q(\abs_multiplicand[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2349_ (.CLK(net1),
    .D(_0045_),
    .Q(\abs_multiplicand[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2350_ (.CLK(net1),
    .D(_0046_),
    .Q(\abs_multiplicand[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2351_ (.CLK(net1),
    .D(_0047_),
    .Q(\abs_multiplicand[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2352_ (.CLK(net1),
    .D(_0048_),
    .Q(\abs_multiplicand[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2353_ (.CLK(net1),
    .D(_0049_),
    .Q(\abs_multiplicand[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2354_ (.CLK(net1),
    .D(_0050_),
    .Q(\abs_multiplicand[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2355_ (.CLK(net1),
    .D(_0051_),
    .Q(\abs_multiplicand[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2356_ (.CLK(net1),
    .D(_0052_),
    .Q(\abs_multiplicand[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2357_ (.CLK(net1),
    .D(_0053_),
    .Q(\abs_multiplicand[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2358_ (.CLK(net1),
    .D(_0054_),
    .Q(\abs_multiplicand[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2359_ (.CLK(net1),
    .D(_0055_),
    .Q(\abs_multiplicand[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2360_ (.CLK(net1),
    .D(_0056_),
    .Q(\abs_multiplicand[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2361_ (.CLK(net1),
    .D(_0057_),
    .Q(\abs_multiplicand[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2362_ (.CLK(net1),
    .D(_0058_),
    .Q(\abs_multiplicand[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2363_ (.CLK(net1),
    .D(_0059_),
    .Q(\abs_multiplicand[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2364_ (.CLK(net1),
    .D(_0060_),
    .Q(\abs_multiplicand[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2365_ (.CLK(net1),
    .D(_0061_),
    .Q(\abs_multiplicand[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2366_ (.CLK(net1),
    .D(_0062_),
    .Q(\abs_multiplicand[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2367_ (.CLK(net1),
    .D(_0063_),
    .Q(\M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2368_ (.CLK(net1),
    .D(_0064_),
    .Q(\M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2369_ (.CLK(net1),
    .D(_0065_),
    .Q(\M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2370_ (.CLK(net1),
    .D(_0066_),
    .Q(\M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2371_ (.CLK(net1),
    .D(_0067_),
    .Q(\M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2372_ (.CLK(net1),
    .D(_0068_),
    .Q(\M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2373_ (.CLK(net1),
    .D(_0069_),
    .Q(\M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2374_ (.CLK(net1),
    .D(_0070_),
    .Q(\M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2375_ (.CLK(net1),
    .D(_0071_),
    .Q(\M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2376_ (.CLK(net1),
    .D(_0072_),
    .Q(\M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2377_ (.CLK(net1),
    .D(_0073_),
    .Q(\M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2378_ (.CLK(net1),
    .D(_0074_),
    .Q(\M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2379_ (.CLK(net1),
    .D(_0075_),
    .Q(\M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2380_ (.CLK(net1),
    .D(_0076_),
    .Q(\M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2381_ (.CLK(net1),
    .D(_0077_),
    .Q(\M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2382_ (.CLK(net1),
    .D(_0078_),
    .Q(\M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2383_ (.CLK(net1),
    .D(_0079_),
    .Q(\M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2384_ (.CLK(net1),
    .D(_0080_),
    .Q(\M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2385_ (.CLK(net1),
    .D(_0081_),
    .Q(\M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2386_ (.CLK(net1),
    .D(_0082_),
    .Q(\M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2387_ (.CLK(net1),
    .D(_0083_),
    .Q(\M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2388_ (.CLK(net1),
    .D(_0084_),
    .Q(\M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2389_ (.CLK(net1),
    .D(_0085_),
    .Q(\M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2390_ (.CLK(net1),
    .D(_0086_),
    .Q(\M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2391_ (.CLK(net1),
    .D(_0087_),
    .Q(\M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2392_ (.CLK(net1),
    .D(_0088_),
    .Q(\M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2393_ (.CLK(net1),
    .D(_0089_),
    .Q(\M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2394_ (.CLK(net1),
    .D(_0090_),
    .Q(\M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2395_ (.CLK(net1),
    .D(_0091_),
    .Q(\M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2396_ (.CLK(net1),
    .D(_0092_),
    .Q(\M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2397_ (.CLK(net1),
    .D(_0093_),
    .Q(\M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2398_ (.CLK(net1),
    .D(_0094_),
    .Q(\M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2399_ (.CLK(net1),
    .D(_0095_),
    .Q(\Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2400_ (.CLK(net1),
    .D(_0096_),
    .Q(\Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2401_ (.CLK(net1),
    .D(_0097_),
    .Q(\Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2402_ (.CLK(net1),
    .D(_0098_),
    .Q(\Q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2403_ (.CLK(net1),
    .D(_0099_),
    .Q(\Q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2404_ (.CLK(net1),
    .D(_0100_),
    .Q(\Q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2405_ (.CLK(net1),
    .D(_0101_),
    .Q(\Q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2406_ (.CLK(net1),
    .D(_0102_),
    .Q(\Q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2407_ (.CLK(net1),
    .D(_0103_),
    .Q(\Q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2408_ (.CLK(net1),
    .D(_0104_),
    .Q(\Q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2409_ (.CLK(net1),
    .D(_0105_),
    .Q(\Q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2410_ (.CLK(net1),
    .D(_0106_),
    .Q(\Q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2411_ (.CLK(net1),
    .D(_0107_),
    .Q(\Q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2412_ (.CLK(net1),
    .D(_0108_),
    .Q(\Q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2413_ (.CLK(net1),
    .D(_0109_),
    .Q(\Q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2414_ (.CLK(net1),
    .D(_0110_),
    .Q(\Q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2415_ (.CLK(net1),
    .D(_0111_),
    .Q(\Q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2416_ (.CLK(net1),
    .D(_0112_),
    .Q(\Q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2417_ (.CLK(net1),
    .D(_0113_),
    .Q(\Q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2418_ (.CLK(net1),
    .D(_0114_),
    .Q(\Q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2419_ (.CLK(net1),
    .D(_0115_),
    .Q(\Q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2420_ (.CLK(net1),
    .D(_0116_),
    .Q(\Q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2421_ (.CLK(net1),
    .D(_0117_),
    .Q(\Q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2422_ (.CLK(net1),
    .D(_0118_),
    .Q(\Q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2423_ (.CLK(net1),
    .D(_0119_),
    .Q(\Q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2424_ (.CLK(net1),
    .D(_0120_),
    .Q(\Q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2425_ (.CLK(net1),
    .D(_0121_),
    .Q(\Q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2426_ (.CLK(net1),
    .D(_0122_),
    .Q(\Q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2427_ (.CLK(net1),
    .D(_0123_),
    .Q(\Q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2428_ (.CLK(net1),
    .D(_0124_),
    .Q(\Q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2429_ (.CLK(net1),
    .D(_0125_),
    .Q(\Q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2430_ (.CLK(net1),
    .D(_0126_),
    .Q(\Q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2431_ (.CLK(net1),
    .D(_0127_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _2432_ (.CLK(net1),
    .D(_0128_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _2433_ (.CLK(net1),
    .D(_0129_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_1 _2434_ (.CLK(net1),
    .D(_0130_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _2435_ (.CLK(net1),
    .D(_0131_),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_1 _2436_ (.CLK(net1),
    .D(_0132_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_1 _2437_ (.CLK(net1),
    .D(_0133_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_1 _2438_ (.CLK(net1),
    .D(_0134_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_1 _2439_ (.CLK(net1),
    .D(_0135_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _2440_ (.CLK(net1),
    .D(_0136_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_1 _2441_ (.CLK(net1),
    .D(_0137_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _2442_ (.CLK(net1),
    .D(_0138_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _2443_ (.CLK(net1),
    .D(_0139_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _2444_ (.CLK(net1),
    .D(_0140_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _2445_ (.CLK(net1),
    .D(_0141_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _2446_ (.CLK(net1),
    .D(_0142_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _2447_ (.CLK(net1),
    .D(_0143_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _2448_ (.CLK(net1),
    .D(_0144_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _2449_ (.CLK(net1),
    .D(_0145_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _2450_ (.CLK(net1),
    .D(_0146_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _2451_ (.CLK(net1),
    .D(_0147_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_1 _2452_ (.CLK(net1),
    .D(_0148_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _2453_ (.CLK(net1),
    .D(_0149_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _2454_ (.CLK(net1),
    .D(_0150_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _2455_ (.CLK(net1),
    .D(_0151_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_1 _2456_ (.CLK(net1),
    .D(_0152_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _2457_ (.CLK(net1),
    .D(_0153_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _2458_ (.CLK(net1),
    .D(_0154_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_1 _2459_ (.CLK(net1),
    .D(_0155_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _2460_ (.CLK(net1),
    .D(_0156_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _2461_ (.CLK(net1),
    .D(_0157_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _2462_ (.CLK(net1),
    .D(_0158_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_1 _2463_ (.CLK(net1),
    .D(_0159_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _2464_ (.CLK(net1),
    .D(_0160_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _2465_ (.CLK(net1),
    .D(_0161_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _2466_ (.CLK(net1),
    .D(_0162_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _2467_ (.CLK(net1),
    .D(_0163_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _2468_ (.CLK(net1),
    .D(_0164_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _2469_ (.CLK(net1),
    .D(_0165_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _2470_ (.CLK(net1),
    .D(_0166_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _2471_ (.CLK(net1),
    .D(_0167_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_1 _2472_ (.CLK(net1),
    .D(_0168_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_1 _2473_ (.CLK(net1),
    .D(_0169_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_1 _2474_ (.CLK(net1),
    .D(_0170_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_1 _2475_ (.CLK(net1),
    .D(_0171_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_1 _2476_ (.CLK(net1),
    .D(_0172_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_1 _2477_ (.CLK(net1),
    .D(_0173_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_1 _2478_ (.CLK(net1),
    .D(_0174_),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_1 _2479_ (.CLK(net1),
    .D(_0175_),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_1 _2480_ (.CLK(net1),
    .D(_0176_),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_1 _2481_ (.CLK(net1),
    .D(_0177_),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_1 _2482_ (.CLK(net1),
    .D(_0178_),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_1 _2483_ (.CLK(net1),
    .D(_0179_),
    .Q(net115));
 sky130_fd_sc_hd__dfxtp_1 _2484_ (.CLK(net1),
    .D(_0180_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_1 _2485_ (.CLK(net1),
    .D(_0181_),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_1 _2486_ (.CLK(net1),
    .D(_0182_),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_1 _2487_ (.CLK(net1),
    .D(_0183_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_1 _2488_ (.CLK(net1),
    .D(_0184_),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_1 _2489_ (.CLK(net1),
    .D(_0185_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_1 _2490_ (.CLK(net1),
    .D(_0186_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_1 _2491_ (.CLK(net1),
    .D(_0187_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_1 _2492_ (.CLK(net1),
    .D(_0188_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_1 _2493_ (.CLK(net1),
    .D(_0189_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_1 _2494_ (.CLK(net1),
    .D(_0190_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_1 _2495_ (.CLK(net1),
    .D(_0191_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _2496_ (.CLK(net1),
    .D(_0192_),
    .Q(\abs_multiplicand[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2497_ (.CLK(net1),
    .D(_0193_),
    .Q(\abs_multiplier[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2498_ (.CLK(net1),
    .D(_0194_),
    .Q(\count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2499_ (.CLK(net1),
    .D(_0195_),
    .Q(\count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2500_ (.CLK(net1),
    .D(_0196_),
    .Q(\count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2501_ (.CLK(net1),
    .D(_0197_),
    .Q(\count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2502_ (.CLK(net1),
    .D(_0198_),
    .Q(\count[4] ));
 sky130_fd_sc_hd__dfxtp_4 _2503_ (.CLK(net1),
    .D(_0199_),
    .Q(\count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2504_ (.CLK(net1),
    .D(_0200_),
    .Q(\A[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2505_ (.CLK(net1),
    .D(_0201_),
    .Q(\A[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2506_ (.CLK(net1),
    .D(_0202_),
    .Q(\A[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2507_ (.CLK(net1),
    .D(_0203_),
    .Q(\A[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2508_ (.CLK(net1),
    .D(_0204_),
    .Q(\A[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2509_ (.CLK(net1),
    .D(_0205_),
    .Q(\A[5] ));
 sky130_fd_sc_hd__dfxtp_2 _2510_ (.CLK(net1),
    .D(_0206_),
    .Q(\A[6] ));
 sky130_fd_sc_hd__dfxtp_2 _2511_ (.CLK(net1),
    .D(_0207_),
    .Q(\A[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2512_ (.CLK(net1),
    .D(_0208_),
    .Q(\A[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2513_ (.CLK(net1),
    .D(_0209_),
    .Q(\A[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2514_ (.CLK(net1),
    .D(_0210_),
    .Q(\A[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2515_ (.CLK(net1),
    .D(_0211_),
    .Q(\A[11] ));
 sky130_fd_sc_hd__dfxtp_2 _2516_ (.CLK(net1),
    .D(_0212_),
    .Q(\A[12] ));
 sky130_fd_sc_hd__dfxtp_2 _2517_ (.CLK(net1),
    .D(_0213_),
    .Q(\A[13] ));
 sky130_fd_sc_hd__dfxtp_2 _2518_ (.CLK(net1),
    .D(_0214_),
    .Q(\A[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2519_ (.CLK(net1),
    .D(_0215_),
    .Q(\A[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2520_ (.CLK(net1),
    .D(_0216_),
    .Q(\A[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2521_ (.CLK(net1),
    .D(_0217_),
    .Q(\A[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2522_ (.CLK(net1),
    .D(_0218_),
    .Q(\A[18] ));
 sky130_fd_sc_hd__dfxtp_2 _2523_ (.CLK(net1),
    .D(_0219_),
    .Q(\A[19] ));
 sky130_fd_sc_hd__dfxtp_2 _2524_ (.CLK(net1),
    .D(_0220_),
    .Q(\A[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2525_ (.CLK(net1),
    .D(_0221_),
    .Q(\A[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2526_ (.CLK(net1),
    .D(_0222_),
    .Q(\A[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2527_ (.CLK(net1),
    .D(_0223_),
    .Q(\A[23] ));
 sky130_fd_sc_hd__dfxtp_2 _2528_ (.CLK(net1),
    .D(_0224_),
    .Q(\A[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2529_ (.CLK(net1),
    .D(_0225_),
    .Q(\A[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2530_ (.CLK(net1),
    .D(_0226_),
    .Q(\A[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2531_ (.CLK(net1),
    .D(_0227_),
    .Q(\A[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2532_ (.CLK(net1),
    .D(_0228_),
    .Q(\A[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2533_ (.CLK(net1),
    .D(_0229_),
    .Q(\A[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2534_ (.CLK(net1),
    .D(_0230_),
    .Q(\A[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2535_ (.CLK(net1),
    .D(_0231_),
    .Q(\A[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2536_ (.CLK(net1),
    .D(_0232_),
    .Q(\A[32] ));
 sky130_fd_sc_hd__dfxtp_1 _2537_ (.CLK(net1),
    .D(_0233_),
    .Q(\A[33] ));
 sky130_fd_sc_hd__dfxtp_1 _2538_ (.CLK(net1),
    .D(_0234_),
    .Q(\A[34] ));
 sky130_fd_sc_hd__dfxtp_1 _2539_ (.CLK(net1),
    .D(_0235_),
    .Q(\A[35] ));
 sky130_fd_sc_hd__dfxtp_1 _2540_ (.CLK(net1),
    .D(_0236_),
    .Q(\A[36] ));
 sky130_fd_sc_hd__dfxtp_1 _2541_ (.CLK(net1),
    .D(_0237_),
    .Q(\A[37] ));
 sky130_fd_sc_hd__dfxtp_1 _2542_ (.CLK(net1),
    .D(_0238_),
    .Q(\A[38] ));
 sky130_fd_sc_hd__dfxtp_1 _2543_ (.CLK(net1),
    .D(_0239_),
    .Q(\A[39] ));
 sky130_fd_sc_hd__dfxtp_1 _2544_ (.CLK(net1),
    .D(_0240_),
    .Q(\A[40] ));
 sky130_fd_sc_hd__dfxtp_1 _2545_ (.CLK(net1),
    .D(_0241_),
    .Q(\A[41] ));
 sky130_fd_sc_hd__dfxtp_1 _2546_ (.CLK(net1),
    .D(_0242_),
    .Q(\A[42] ));
 sky130_fd_sc_hd__dfxtp_1 _2547_ (.CLK(net1),
    .D(_0243_),
    .Q(\A[43] ));
 sky130_fd_sc_hd__dfxtp_1 _2548_ (.CLK(net1),
    .D(_0244_),
    .Q(\A[44] ));
 sky130_fd_sc_hd__dfxtp_1 _2549_ (.CLK(net1),
    .D(_0245_),
    .Q(\A[45] ));
 sky130_fd_sc_hd__dfxtp_1 _2550_ (.CLK(net1),
    .D(_0246_),
    .Q(\A[46] ));
 sky130_fd_sc_hd__dfxtp_1 _2551_ (.CLK(net1),
    .D(_0247_),
    .Q(\A[47] ));
 sky130_fd_sc_hd__dfxtp_1 _2552_ (.CLK(net1),
    .D(_0248_),
    .Q(\A[48] ));
 sky130_fd_sc_hd__dfxtp_1 _2553_ (.CLK(net1),
    .D(_0249_),
    .Q(\A[49] ));
 sky130_fd_sc_hd__dfxtp_1 _2554_ (.CLK(net1),
    .D(_0250_),
    .Q(\A[50] ));
 sky130_fd_sc_hd__dfxtp_1 _2555_ (.CLK(net1),
    .D(_0251_),
    .Q(\A[51] ));
 sky130_fd_sc_hd__dfxtp_1 _2556_ (.CLK(net1),
    .D(_0252_),
    .Q(\A[52] ));
 sky130_fd_sc_hd__dfxtp_1 _2557_ (.CLK(net1),
    .D(_0253_),
    .Q(\A[53] ));
 sky130_fd_sc_hd__dfxtp_1 _2558_ (.CLK(net1),
    .D(_0254_),
    .Q(\A[54] ));
 sky130_fd_sc_hd__dfxtp_1 _2559_ (.CLK(net1),
    .D(_0255_),
    .Q(\A[55] ));
 sky130_fd_sc_hd__dfxtp_1 _2560_ (.CLK(net1),
    .D(_0256_),
    .Q(\A[56] ));
 sky130_fd_sc_hd__dfxtp_1 _2561_ (.CLK(net1),
    .D(_0257_),
    .Q(\A[57] ));
 sky130_fd_sc_hd__dfxtp_1 _2562_ (.CLK(net1),
    .D(_0258_),
    .Q(\A[58] ));
 sky130_fd_sc_hd__dfxtp_1 _2563_ (.CLK(net1),
    .D(_0259_),
    .Q(\A[59] ));
 sky130_fd_sc_hd__dfxtp_1 _2564_ (.CLK(net1),
    .D(_0260_),
    .Q(\A[60] ));
 sky130_fd_sc_hd__dfxtp_1 _2565_ (.CLK(net1),
    .D(_0261_),
    .Q(\A[61] ));
 sky130_fd_sc_hd__dfxtp_1 _2566_ (.CLK(net1),
    .D(_0262_),
    .Q(\A[62] ));
 sky130_fd_sc_hd__clkbuf_16 input1 (.A(clk),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(multiplicand[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(multiplicand[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(multiplicand[11]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(multiplicand[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(multiplicand[13]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(multiplicand[14]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(multiplicand[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(multiplicand[16]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(multiplicand[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(multiplicand[18]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(multiplicand[19]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(multiplicand[1]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(multiplicand[20]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(multiplicand[21]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(multiplicand[22]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(multiplicand[23]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(multiplicand[24]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(multiplicand[25]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(multiplicand[26]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(multiplicand[27]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(multiplicand[28]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(multiplicand[29]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(multiplicand[2]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(multiplicand[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_16 input26 (.A(multiplicand[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(multiplicand[3]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(multiplicand[4]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(multiplicand[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(multiplicand[6]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(multiplicand[7]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(multiplicand[8]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(multiplicand[9]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(multiplier[0]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(multiplier[10]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(multiplier[11]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(multiplier[12]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(multiplier[13]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(multiplier[14]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(multiplier[15]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(multiplier[16]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(multiplier[17]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(multiplier[18]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(multiplier[19]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(multiplier[1]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(multiplier[20]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(multiplier[21]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(multiplier[22]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(multiplier[23]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(multiplier[24]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(multiplier[25]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(multiplier[26]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(multiplier[27]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(multiplier[28]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(multiplier[29]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(multiplier[2]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(multiplier[30]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_16 input58 (.A(multiplier[31]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(multiplier[3]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(multiplier[4]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(multiplier[5]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(multiplier[6]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(multiplier[7]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(multiplier[8]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(multiplier[9]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_16 input66 (.A(rst),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_16 output67 (.A(net67),
    .X(done));
 sky130_fd_sc_hd__clkbuf_16 output68 (.A(net68),
    .X(product[0]));
 sky130_fd_sc_hd__clkbuf_16 output69 (.A(net69),
    .X(product[10]));
 sky130_fd_sc_hd__clkbuf_16 output70 (.A(net70),
    .X(product[11]));
 sky130_fd_sc_hd__clkbuf_16 output71 (.A(net71),
    .X(product[12]));
 sky130_fd_sc_hd__clkbuf_16 output72 (.A(net72),
    .X(product[13]));
 sky130_fd_sc_hd__clkbuf_16 output73 (.A(net73),
    .X(product[14]));
 sky130_fd_sc_hd__clkbuf_16 output74 (.A(net74),
    .X(product[15]));
 sky130_fd_sc_hd__clkbuf_16 output75 (.A(net75),
    .X(product[16]));
 sky130_fd_sc_hd__clkbuf_16 output76 (.A(net76),
    .X(product[17]));
 sky130_fd_sc_hd__clkbuf_16 output77 (.A(net77),
    .X(product[18]));
 sky130_fd_sc_hd__clkbuf_16 output78 (.A(net78),
    .X(product[19]));
 sky130_fd_sc_hd__clkbuf_16 output79 (.A(net79),
    .X(product[1]));
 sky130_fd_sc_hd__clkbuf_16 output80 (.A(net80),
    .X(product[20]));
 sky130_fd_sc_hd__clkbuf_16 output81 (.A(net81),
    .X(product[21]));
 sky130_fd_sc_hd__clkbuf_16 output82 (.A(net82),
    .X(product[22]));
 sky130_fd_sc_hd__clkbuf_16 output83 (.A(net83),
    .X(product[23]));
 sky130_fd_sc_hd__clkbuf_16 output84 (.A(net84),
    .X(product[24]));
 sky130_fd_sc_hd__clkbuf_16 output85 (.A(net85),
    .X(product[25]));
 sky130_fd_sc_hd__clkbuf_16 output86 (.A(net86),
    .X(product[26]));
 sky130_fd_sc_hd__clkbuf_16 output87 (.A(net87),
    .X(product[27]));
 sky130_fd_sc_hd__clkbuf_16 output88 (.A(net88),
    .X(product[28]));
 sky130_fd_sc_hd__clkbuf_16 output89 (.A(net89),
    .X(product[29]));
 sky130_fd_sc_hd__clkbuf_16 output90 (.A(net90),
    .X(product[2]));
 sky130_fd_sc_hd__clkbuf_16 output91 (.A(net91),
    .X(product[30]));
 sky130_fd_sc_hd__clkbuf_16 output92 (.A(net92),
    .X(product[31]));
 sky130_fd_sc_hd__clkbuf_16 output93 (.A(net93),
    .X(product[32]));
 sky130_fd_sc_hd__clkbuf_16 output94 (.A(net94),
    .X(product[33]));
 sky130_fd_sc_hd__clkbuf_16 output95 (.A(net95),
    .X(product[34]));
 sky130_fd_sc_hd__clkbuf_16 output96 (.A(net96),
    .X(product[35]));
 sky130_fd_sc_hd__clkbuf_16 output97 (.A(net97),
    .X(product[36]));
 sky130_fd_sc_hd__clkbuf_16 output98 (.A(net98),
    .X(product[37]));
 sky130_fd_sc_hd__clkbuf_16 output99 (.A(net99),
    .X(product[38]));
 sky130_fd_sc_hd__clkbuf_16 output100 (.A(net100),
    .X(product[39]));
 sky130_fd_sc_hd__clkbuf_16 output101 (.A(net101),
    .X(product[3]));
 sky130_fd_sc_hd__clkbuf_16 output102 (.A(net102),
    .X(product[40]));
 sky130_fd_sc_hd__clkbuf_16 output103 (.A(net103),
    .X(product[41]));
 sky130_fd_sc_hd__clkbuf_16 output104 (.A(net104),
    .X(product[42]));
 sky130_fd_sc_hd__clkbuf_16 output105 (.A(net105),
    .X(product[43]));
 sky130_fd_sc_hd__clkbuf_16 output106 (.A(net106),
    .X(product[44]));
 sky130_fd_sc_hd__clkbuf_16 output107 (.A(net107),
    .X(product[45]));
 sky130_fd_sc_hd__clkbuf_16 output108 (.A(net108),
    .X(product[46]));
 sky130_fd_sc_hd__clkbuf_16 output109 (.A(net109),
    .X(product[47]));
 sky130_fd_sc_hd__clkbuf_16 output110 (.A(net110),
    .X(product[48]));
 sky130_fd_sc_hd__clkbuf_16 output111 (.A(net111),
    .X(product[49]));
 sky130_fd_sc_hd__clkbuf_16 output112 (.A(net112),
    .X(product[4]));
 sky130_fd_sc_hd__clkbuf_16 output113 (.A(net113),
    .X(product[50]));
 sky130_fd_sc_hd__clkbuf_16 output114 (.A(net114),
    .X(product[51]));
 sky130_fd_sc_hd__clkbuf_16 output115 (.A(net115),
    .X(product[52]));
 sky130_fd_sc_hd__clkbuf_16 output116 (.A(net116),
    .X(product[53]));
 sky130_fd_sc_hd__clkbuf_16 output117 (.A(net117),
    .X(product[54]));
 sky130_fd_sc_hd__clkbuf_16 output118 (.A(net118),
    .X(product[55]));
 sky130_fd_sc_hd__clkbuf_16 output119 (.A(net119),
    .X(product[56]));
 sky130_fd_sc_hd__clkbuf_16 output120 (.A(net120),
    .X(product[57]));
 sky130_fd_sc_hd__clkbuf_16 output121 (.A(net121),
    .X(product[58]));
 sky130_fd_sc_hd__clkbuf_16 output122 (.A(net122),
    .X(product[59]));
 sky130_fd_sc_hd__clkbuf_16 output123 (.A(net123),
    .X(product[5]));
 sky130_fd_sc_hd__clkbuf_16 output124 (.A(net124),
    .X(product[60]));
 sky130_fd_sc_hd__clkbuf_16 output125 (.A(net125),
    .X(product[61]));
 sky130_fd_sc_hd__clkbuf_16 output126 (.A(net126),
    .X(product[62]));
 sky130_fd_sc_hd__clkbuf_16 output127 (.A(net127),
    .X(product[63]));
 sky130_fd_sc_hd__clkbuf_16 output128 (.A(net128),
    .X(product[6]));
 sky130_fd_sc_hd__clkbuf_16 output129 (.A(net129),
    .X(product[7]));
 sky130_fd_sc_hd__clkbuf_16 output130 (.A(net130),
    .X(product[8]));
 sky130_fd_sc_hd__clkbuf_16 output131 (.A(net131),
    .X(product[9]));
 sky130_fd_sc_hd__buf_12 max_cap132 (.A(_1149_),
    .X(net132));
 sky130_fd_sc_hd__buf_12 max_cap133 (.A(_1049_),
    .X(net133));
 sky130_fd_sc_hd__buf_12 max_cap134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_12 max_cap135 (.A(\count[5] ),
    .X(net135));
endmodule
